##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar  7 18:05:08 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_160b_w16
  CLASS BLOCK ;
  SIZE 243.0000 BY 241.4000 ;
  FOREIGN sram_160b_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 118.1500 0.6000 118.2500 ;
    END
  END CLK
  PIN D[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.6500 0.0000 57.7500 0.6000 ;
    END
  END D[159]
  PIN D[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.4500 0.0000 58.5500 0.6000 ;
    END
  END D[158]
  PIN D[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 59.2500 0.0000 59.3500 0.6000 ;
    END
  END D[157]
  PIN D[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.0500 0.0000 60.1500 0.6000 ;
    END
  END D[156]
  PIN D[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.8500 0.0000 60.9500 0.6000 ;
    END
  END D[155]
  PIN D[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.6500 0.0000 61.7500 0.6000 ;
    END
  END D[154]
  PIN D[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 62.4500 0.0000 62.5500 0.6000 ;
    END
  END D[153]
  PIN D[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.2500 0.0000 63.3500 0.6000 ;
    END
  END D[152]
  PIN D[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64.0500 0.0000 64.1500 0.6000 ;
    END
  END D[151]
  PIN D[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64.8500 0.0000 64.9500 0.6000 ;
    END
  END D[150]
  PIN D[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.6500 0.0000 65.7500 0.6000 ;
    END
  END D[149]
  PIN D[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.4500 0.0000 66.5500 0.6000 ;
    END
  END D[148]
  PIN D[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 67.2500 0.0000 67.3500 0.6000 ;
    END
  END D[147]
  PIN D[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.0500 0.0000 68.1500 0.6000 ;
    END
  END D[146]
  PIN D[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.8500 0.0000 68.9500 0.6000 ;
    END
  END D[145]
  PIN D[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.6500 0.0000 69.7500 0.6000 ;
    END
  END D[144]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.4500 0.0000 70.5500 0.6000 ;
    END
  END D[143]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.2500 0.0000 71.3500 0.6000 ;
    END
  END D[142]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 72.0500 0.0000 72.1500 0.6000 ;
    END
  END D[141]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 72.8500 0.0000 72.9500 0.6000 ;
    END
  END D[140]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.6500 0.0000 73.7500 0.6000 ;
    END
  END D[139]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.4500 0.0000 74.5500 0.6000 ;
    END
  END D[138]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 75.2500 0.0000 75.3500 0.6000 ;
    END
  END D[137]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.0500 0.0000 76.1500 0.6000 ;
    END
  END D[136]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.8500 0.0000 76.9500 0.6000 ;
    END
  END D[135]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.6500 0.0000 77.7500 0.6000 ;
    END
  END D[134]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 78.4500 0.0000 78.5500 0.6000 ;
    END
  END D[133]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.2500 0.0000 79.3500 0.6000 ;
    END
  END D[132]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.0500 0.0000 80.1500 0.6000 ;
    END
  END D[131]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.8500 0.0000 80.9500 0.6000 ;
    END
  END D[130]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.6500 0.0000 81.7500 0.6000 ;
    END
  END D[129]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.4500 0.0000 82.5500 0.6000 ;
    END
  END D[128]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 83.2500 0.0000 83.3500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.0500 0.0000 84.1500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.8500 0.0000 84.9500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.6500 0.0000 85.7500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.4500 0.0000 86.5500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.2500 0.0000 87.3500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.0500 0.0000 88.1500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.8500 0.0000 88.9500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.6500 0.0000 89.7500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.4500 0.0000 90.5500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.2500 0.0000 91.3500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.0500 0.0000 92.1500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.8500 0.0000 92.9500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.6500 0.0000 93.7500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 94.4500 0.0000 94.5500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.2500 0.0000 95.3500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.0500 0.0000 96.1500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.8500 0.0000 96.9500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.6500 0.0000 97.7500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.4500 0.0000 98.5500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 99.2500 0.0000 99.3500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.0500 0.0000 100.1500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.8500 0.0000 100.9500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.6500 0.0000 101.7500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 102.4500 0.0000 102.5500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.2500 0.0000 103.3500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.0500 0.0000 104.1500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.8500 0.0000 104.9500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.6500 0.0000 105.7500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.4500 0.0000 106.5500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 107.2500 0.0000 107.3500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.0500 0.0000 108.1500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.8500 0.0000 108.9500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.6500 0.0000 109.7500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 110.4500 0.0000 110.5500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.2500 0.0000 111.3500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.0500 0.0000 112.1500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.8500 0.0000 112.9500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.6500 0.0000 113.7500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.4500 0.0000 114.5500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.2500 0.0000 115.3500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.0500 0.0000 116.1500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.8500 0.0000 116.9500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.6500 0.0000 117.7500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 118.4500 0.0000 118.5500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.2500 0.0000 119.3500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.0500 0.0000 120.1500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.8500 0.0000 120.9500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.6500 0.0000 121.7500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.4500 0.0000 122.5500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.2500 0.0000 123.3500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.0500 0.0000 124.1500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.8500 0.0000 124.9500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.6500 0.0000 125.7500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 126.4500 0.0000 126.5500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.2500 0.0000 127.3500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.0500 0.0000 128.1500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.8500 0.0000 128.9500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.6500 0.0000 129.7500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.4500 0.0000 130.5500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.2500 0.0000 131.3500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.0500 0.0000 132.1500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.8500 0.0000 132.9500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.6500 0.0000 133.7500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.4500 0.0000 134.5500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.2500 0.0000 135.3500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.0500 0.0000 136.1500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.8500 0.0000 136.9500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.6500 0.0000 137.7500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.4500 0.0000 138.5500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 139.2500 0.0000 139.3500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.0500 0.0000 140.1500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.8500 0.0000 140.9500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.6500 0.0000 141.7500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 142.4500 0.0000 142.5500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.2500 0.0000 143.3500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.0500 0.0000 144.1500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.8500 0.0000 144.9500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.6500 0.0000 145.7500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.4500 0.0000 146.5500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.2500 0.0000 147.3500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.0500 0.0000 148.1500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.8500 0.0000 148.9500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.6500 0.0000 149.7500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.4500 0.0000 150.5500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.2500 0.0000 151.3500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.0500 0.0000 152.1500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.8500 0.0000 152.9500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.6500 0.0000 153.7500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.4500 0.0000 154.5500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.2500 0.0000 155.3500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.0500 0.0000 156.1500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.8500 0.0000 156.9500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.6500 0.0000 157.7500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.4500 0.0000 158.5500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.2500 0.0000 159.3500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.0500 0.0000 160.1500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.8500 0.0000 160.9500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.6500 0.0000 161.7500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.4500 0.0000 162.5500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.2500 0.0000 163.3500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.0500 0.0000 164.1500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.8500 0.0000 164.9500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.6500 0.0000 165.7500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.4500 0.0000 166.5500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.2500 0.0000 167.3500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.0500 0.0000 168.1500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.8500 0.0000 168.9500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.6500 0.0000 169.7500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.4500 0.0000 170.5500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.2500 0.0000 171.3500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.0500 0.0000 172.1500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.8500 0.0000 172.9500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.6500 0.0000 173.7500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.4500 0.0000 174.5500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.2500 0.0000 175.3500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.0500 0.0000 176.1500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.8500 0.0000 176.9500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.6500 0.0000 177.7500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.4500 0.0000 178.5500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.2500 0.0000 179.3500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.0500 0.0000 180.1500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.8500 0.0000 180.9500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.6500 0.0000 181.7500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.4500 0.0000 182.5500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.2500 0.0000 183.3500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.0500 0.0000 184.1500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.8500 0.0000 184.9500 0.6000 ;
    END
  END D[0]
  PIN Q[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 57.6500 240.8000 57.7500 241.4000 ;
    END
  END Q[159]
  PIN Q[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 58.4500 240.8000 58.5500 241.4000 ;
    END
  END Q[158]
  PIN Q[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 59.2500 240.8000 59.3500 241.4000 ;
    END
  END Q[157]
  PIN Q[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.0500 240.8000 60.1500 241.4000 ;
    END
  END Q[156]
  PIN Q[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 60.8500 240.8000 60.9500 241.4000 ;
    END
  END Q[155]
  PIN Q[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 61.6500 240.8000 61.7500 241.4000 ;
    END
  END Q[154]
  PIN Q[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 62.4500 240.8000 62.5500 241.4000 ;
    END
  END Q[153]
  PIN Q[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 63.2500 240.8000 63.3500 241.4000 ;
    END
  END Q[152]
  PIN Q[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64.0500 240.8000 64.1500 241.4000 ;
    END
  END Q[151]
  PIN Q[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 64.8500 240.8000 64.9500 241.4000 ;
    END
  END Q[150]
  PIN Q[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 65.6500 240.8000 65.7500 241.4000 ;
    END
  END Q[149]
  PIN Q[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.4500 240.8000 66.5500 241.4000 ;
    END
  END Q[148]
  PIN Q[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 67.2500 240.8000 67.3500 241.4000 ;
    END
  END Q[147]
  PIN Q[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.0500 240.8000 68.1500 241.4000 ;
    END
  END Q[146]
  PIN Q[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 68.8500 240.8000 68.9500 241.4000 ;
    END
  END Q[145]
  PIN Q[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.6500 240.8000 69.7500 241.4000 ;
    END
  END Q[144]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.4500 240.8000 70.5500 241.4000 ;
    END
  END Q[143]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.2500 240.8000 71.3500 241.4000 ;
    END
  END Q[142]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 72.0500 240.8000 72.1500 241.4000 ;
    END
  END Q[141]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 72.8500 240.8000 72.9500 241.4000 ;
    END
  END Q[140]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.6500 240.8000 73.7500 241.4000 ;
    END
  END Q[139]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.4500 240.8000 74.5500 241.4000 ;
    END
  END Q[138]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 75.2500 240.8000 75.3500 241.4000 ;
    END
  END Q[137]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.0500 240.8000 76.1500 241.4000 ;
    END
  END Q[136]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.8500 240.8000 76.9500 241.4000 ;
    END
  END Q[135]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.6500 240.8000 77.7500 241.4000 ;
    END
  END Q[134]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 78.4500 240.8000 78.5500 241.4000 ;
    END
  END Q[133]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.2500 240.8000 79.3500 241.4000 ;
    END
  END Q[132]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.0500 240.8000 80.1500 241.4000 ;
    END
  END Q[131]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.8500 240.8000 80.9500 241.4000 ;
    END
  END Q[130]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.6500 240.8000 81.7500 241.4000 ;
    END
  END Q[129]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.4500 240.8000 82.5500 241.4000 ;
    END
  END Q[128]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 83.2500 240.8000 83.3500 241.4000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.0500 240.8000 84.1500 241.4000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.8500 240.8000 84.9500 241.4000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.6500 240.8000 85.7500 241.4000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.4500 240.8000 86.5500 241.4000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.2500 240.8000 87.3500 241.4000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.0500 240.8000 88.1500 241.4000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.8500 240.8000 88.9500 241.4000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.6500 240.8000 89.7500 241.4000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.4500 240.8000 90.5500 241.4000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.2500 240.8000 91.3500 241.4000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.0500 240.8000 92.1500 241.4000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.8500 240.8000 92.9500 241.4000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.6500 240.8000 93.7500 241.4000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 94.4500 240.8000 94.5500 241.4000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.2500 240.8000 95.3500 241.4000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.0500 240.8000 96.1500 241.4000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.8500 240.8000 96.9500 241.4000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.6500 240.8000 97.7500 241.4000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.4500 240.8000 98.5500 241.4000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 99.2500 240.8000 99.3500 241.4000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.0500 240.8000 100.1500 241.4000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.8500 240.8000 100.9500 241.4000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.6500 240.8000 101.7500 241.4000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 102.4500 240.8000 102.5500 241.4000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.2500 240.8000 103.3500 241.4000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.0500 240.8000 104.1500 241.4000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.8500 240.8000 104.9500 241.4000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.6500 240.8000 105.7500 241.4000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.4500 240.8000 106.5500 241.4000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 107.2500 240.8000 107.3500 241.4000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.0500 240.8000 108.1500 241.4000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.8500 240.8000 108.9500 241.4000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.6500 240.8000 109.7500 241.4000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 110.4500 240.8000 110.5500 241.4000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.2500 240.8000 111.3500 241.4000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.0500 240.8000 112.1500 241.4000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.8500 240.8000 112.9500 241.4000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.6500 240.8000 113.7500 241.4000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.4500 240.8000 114.5500 241.4000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.2500 240.8000 115.3500 241.4000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.0500 240.8000 116.1500 241.4000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.8500 240.8000 116.9500 241.4000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.6500 240.8000 117.7500 241.4000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 118.4500 240.8000 118.5500 241.4000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.2500 240.8000 119.3500 241.4000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.0500 240.8000 120.1500 241.4000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.8500 240.8000 120.9500 241.4000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.6500 240.8000 121.7500 241.4000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.4500 240.8000 122.5500 241.4000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.2500 240.8000 123.3500 241.4000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.0500 240.8000 124.1500 241.4000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.8500 240.8000 124.9500 241.4000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.6500 240.8000 125.7500 241.4000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 126.4500 240.8000 126.5500 241.4000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.2500 240.8000 127.3500 241.4000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.0500 240.8000 128.1500 241.4000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.8500 240.8000 128.9500 241.4000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.6500 240.8000 129.7500 241.4000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.4500 240.8000 130.5500 241.4000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.2500 240.8000 131.3500 241.4000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.0500 240.8000 132.1500 241.4000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.8500 240.8000 132.9500 241.4000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.6500 240.8000 133.7500 241.4000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.4500 240.8000 134.5500 241.4000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.2500 240.8000 135.3500 241.4000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.0500 240.8000 136.1500 241.4000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.8500 240.8000 136.9500 241.4000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.6500 240.8000 137.7500 241.4000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.4500 240.8000 138.5500 241.4000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 139.2500 240.8000 139.3500 241.4000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.0500 240.8000 140.1500 241.4000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.8500 240.8000 140.9500 241.4000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.6500 240.8000 141.7500 241.4000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 142.4500 240.8000 142.5500 241.4000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.2500 240.8000 143.3500 241.4000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.0500 240.8000 144.1500 241.4000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.8500 240.8000 144.9500 241.4000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.6500 240.8000 145.7500 241.4000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.4500 240.8000 146.5500 241.4000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.2500 240.8000 147.3500 241.4000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.0500 240.8000 148.1500 241.4000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.8500 240.8000 148.9500 241.4000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.6500 240.8000 149.7500 241.4000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.4500 240.8000 150.5500 241.4000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.2500 240.8000 151.3500 241.4000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.0500 240.8000 152.1500 241.4000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.8500 240.8000 152.9500 241.4000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.6500 240.8000 153.7500 241.4000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.4500 240.8000 154.5500 241.4000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.2500 240.8000 155.3500 241.4000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.0500 240.8000 156.1500 241.4000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.8500 240.8000 156.9500 241.4000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.6500 240.8000 157.7500 241.4000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.4500 240.8000 158.5500 241.4000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.2500 240.8000 159.3500 241.4000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.0500 240.8000 160.1500 241.4000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.8500 240.8000 160.9500 241.4000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.6500 240.8000 161.7500 241.4000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.4500 240.8000 162.5500 241.4000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.2500 240.8000 163.3500 241.4000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.0500 240.8000 164.1500 241.4000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.8500 240.8000 164.9500 241.4000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.6500 240.8000 165.7500 241.4000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.4500 240.8000 166.5500 241.4000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.2500 240.8000 167.3500 241.4000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.0500 240.8000 168.1500 241.4000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.8500 240.8000 168.9500 241.4000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.6500 240.8000 169.7500 241.4000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.4500 240.8000 170.5500 241.4000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.2500 240.8000 171.3500 241.4000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.0500 240.8000 172.1500 241.4000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.8500 240.8000 172.9500 241.4000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.6500 240.8000 173.7500 241.4000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.4500 240.8000 174.5500 241.4000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.2500 240.8000 175.3500 241.4000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.0500 240.8000 176.1500 241.4000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.8500 240.8000 176.9500 241.4000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.6500 240.8000 177.7500 241.4000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.4500 240.8000 178.5500 241.4000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.2500 240.8000 179.3500 241.4000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.0500 240.8000 180.1500 241.4000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.8500 240.8000 180.9500 241.4000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.6500 240.8000 181.7500 241.4000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.4500 240.8000 182.5500 241.4000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.2500 240.8000 183.3500 241.4000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.0500 240.8000 184.1500 241.4000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.8500 240.8000 184.9500 241.4000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 122.1500 0.6000 122.2500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 122.9500 0.6000 123.0500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 118.9500 0.6000 119.0500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 119.7500 0.6000 119.8500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 120.5500 0.6000 120.6500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 121.3500 0.6000 121.4500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 239.0000 1.0000 240.0000 240.4000 ;
        RECT 1.0000 1.0000 2.0000 240.4000 ;
        RECT 1.0000 240.2350 2.0000 240.5650 ;
        RECT 239.0000 240.2350 240.0000 240.5650 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 241.0000 1.0000 242.0000 240.4000 ;
        RECT 3.0000 1.0000 4.0000 240.4000 ;
        RECT 3.0000 0.8350 4.0000 1.1650 ;
        RECT 241.0000 0.8350 242.0000 1.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 243.0000 241.4000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 243.0000 241.4000 ;
    LAYER M3 ;
      RECT 185.1100 240.6400 243.0000 241.4000 ;
      RECT 184.3100 240.6400 184.6900 241.4000 ;
      RECT 183.5100 240.6400 183.8900 241.4000 ;
      RECT 182.7100 240.6400 183.0900 241.4000 ;
      RECT 181.9100 240.6400 182.2900 241.4000 ;
      RECT 181.1100 240.6400 181.4900 241.4000 ;
      RECT 180.3100 240.6400 180.6900 241.4000 ;
      RECT 179.5100 240.6400 179.8900 241.4000 ;
      RECT 178.7100 240.6400 179.0900 241.4000 ;
      RECT 177.9100 240.6400 178.2900 241.4000 ;
      RECT 177.1100 240.6400 177.4900 241.4000 ;
      RECT 176.3100 240.6400 176.6900 241.4000 ;
      RECT 175.5100 240.6400 175.8900 241.4000 ;
      RECT 174.7100 240.6400 175.0900 241.4000 ;
      RECT 173.9100 240.6400 174.2900 241.4000 ;
      RECT 173.1100 240.6400 173.4900 241.4000 ;
      RECT 172.3100 240.6400 172.6900 241.4000 ;
      RECT 171.5100 240.6400 171.8900 241.4000 ;
      RECT 170.7100 240.6400 171.0900 241.4000 ;
      RECT 169.9100 240.6400 170.2900 241.4000 ;
      RECT 169.1100 240.6400 169.4900 241.4000 ;
      RECT 168.3100 240.6400 168.6900 241.4000 ;
      RECT 167.5100 240.6400 167.8900 241.4000 ;
      RECT 166.7100 240.6400 167.0900 241.4000 ;
      RECT 165.9100 240.6400 166.2900 241.4000 ;
      RECT 165.1100 240.6400 165.4900 241.4000 ;
      RECT 164.3100 240.6400 164.6900 241.4000 ;
      RECT 163.5100 240.6400 163.8900 241.4000 ;
      RECT 162.7100 240.6400 163.0900 241.4000 ;
      RECT 161.9100 240.6400 162.2900 241.4000 ;
      RECT 161.1100 240.6400 161.4900 241.4000 ;
      RECT 160.3100 240.6400 160.6900 241.4000 ;
      RECT 159.5100 240.6400 159.8900 241.4000 ;
      RECT 158.7100 240.6400 159.0900 241.4000 ;
      RECT 157.9100 240.6400 158.2900 241.4000 ;
      RECT 157.1100 240.6400 157.4900 241.4000 ;
      RECT 156.3100 240.6400 156.6900 241.4000 ;
      RECT 155.5100 240.6400 155.8900 241.4000 ;
      RECT 154.7100 240.6400 155.0900 241.4000 ;
      RECT 153.9100 240.6400 154.2900 241.4000 ;
      RECT 153.1100 240.6400 153.4900 241.4000 ;
      RECT 152.3100 240.6400 152.6900 241.4000 ;
      RECT 151.5100 240.6400 151.8900 241.4000 ;
      RECT 150.7100 240.6400 151.0900 241.4000 ;
      RECT 149.9100 240.6400 150.2900 241.4000 ;
      RECT 149.1100 240.6400 149.4900 241.4000 ;
      RECT 148.3100 240.6400 148.6900 241.4000 ;
      RECT 147.5100 240.6400 147.8900 241.4000 ;
      RECT 146.7100 240.6400 147.0900 241.4000 ;
      RECT 145.9100 240.6400 146.2900 241.4000 ;
      RECT 145.1100 240.6400 145.4900 241.4000 ;
      RECT 144.3100 240.6400 144.6900 241.4000 ;
      RECT 143.5100 240.6400 143.8900 241.4000 ;
      RECT 142.7100 240.6400 143.0900 241.4000 ;
      RECT 141.9100 240.6400 142.2900 241.4000 ;
      RECT 141.1100 240.6400 141.4900 241.4000 ;
      RECT 140.3100 240.6400 140.6900 241.4000 ;
      RECT 139.5100 240.6400 139.8900 241.4000 ;
      RECT 138.7100 240.6400 139.0900 241.4000 ;
      RECT 137.9100 240.6400 138.2900 241.4000 ;
      RECT 137.1100 240.6400 137.4900 241.4000 ;
      RECT 136.3100 240.6400 136.6900 241.4000 ;
      RECT 135.5100 240.6400 135.8900 241.4000 ;
      RECT 134.7100 240.6400 135.0900 241.4000 ;
      RECT 133.9100 240.6400 134.2900 241.4000 ;
      RECT 133.1100 240.6400 133.4900 241.4000 ;
      RECT 132.3100 240.6400 132.6900 241.4000 ;
      RECT 131.5100 240.6400 131.8900 241.4000 ;
      RECT 130.7100 240.6400 131.0900 241.4000 ;
      RECT 129.9100 240.6400 130.2900 241.4000 ;
      RECT 129.1100 240.6400 129.4900 241.4000 ;
      RECT 128.3100 240.6400 128.6900 241.4000 ;
      RECT 127.5100 240.6400 127.8900 241.4000 ;
      RECT 126.7100 240.6400 127.0900 241.4000 ;
      RECT 125.9100 240.6400 126.2900 241.4000 ;
      RECT 125.1100 240.6400 125.4900 241.4000 ;
      RECT 124.3100 240.6400 124.6900 241.4000 ;
      RECT 123.5100 240.6400 123.8900 241.4000 ;
      RECT 122.7100 240.6400 123.0900 241.4000 ;
      RECT 121.9100 240.6400 122.2900 241.4000 ;
      RECT 121.1100 240.6400 121.4900 241.4000 ;
      RECT 120.3100 240.6400 120.6900 241.4000 ;
      RECT 119.5100 240.6400 119.8900 241.4000 ;
      RECT 118.7100 240.6400 119.0900 241.4000 ;
      RECT 117.9100 240.6400 118.2900 241.4000 ;
      RECT 117.1100 240.6400 117.4900 241.4000 ;
      RECT 116.3100 240.6400 116.6900 241.4000 ;
      RECT 115.5100 240.6400 115.8900 241.4000 ;
      RECT 114.7100 240.6400 115.0900 241.4000 ;
      RECT 113.9100 240.6400 114.2900 241.4000 ;
      RECT 113.1100 240.6400 113.4900 241.4000 ;
      RECT 112.3100 240.6400 112.6900 241.4000 ;
      RECT 111.5100 240.6400 111.8900 241.4000 ;
      RECT 110.7100 240.6400 111.0900 241.4000 ;
      RECT 109.9100 240.6400 110.2900 241.4000 ;
      RECT 109.1100 240.6400 109.4900 241.4000 ;
      RECT 108.3100 240.6400 108.6900 241.4000 ;
      RECT 107.5100 240.6400 107.8900 241.4000 ;
      RECT 106.7100 240.6400 107.0900 241.4000 ;
      RECT 105.9100 240.6400 106.2900 241.4000 ;
      RECT 105.1100 240.6400 105.4900 241.4000 ;
      RECT 104.3100 240.6400 104.6900 241.4000 ;
      RECT 103.5100 240.6400 103.8900 241.4000 ;
      RECT 102.7100 240.6400 103.0900 241.4000 ;
      RECT 101.9100 240.6400 102.2900 241.4000 ;
      RECT 101.1100 240.6400 101.4900 241.4000 ;
      RECT 100.3100 240.6400 100.6900 241.4000 ;
      RECT 99.5100 240.6400 99.8900 241.4000 ;
      RECT 98.7100 240.6400 99.0900 241.4000 ;
      RECT 97.9100 240.6400 98.2900 241.4000 ;
      RECT 97.1100 240.6400 97.4900 241.4000 ;
      RECT 96.3100 240.6400 96.6900 241.4000 ;
      RECT 95.5100 240.6400 95.8900 241.4000 ;
      RECT 94.7100 240.6400 95.0900 241.4000 ;
      RECT 93.9100 240.6400 94.2900 241.4000 ;
      RECT 93.1100 240.6400 93.4900 241.4000 ;
      RECT 92.3100 240.6400 92.6900 241.4000 ;
      RECT 91.5100 240.6400 91.8900 241.4000 ;
      RECT 90.7100 240.6400 91.0900 241.4000 ;
      RECT 89.9100 240.6400 90.2900 241.4000 ;
      RECT 89.1100 240.6400 89.4900 241.4000 ;
      RECT 88.3100 240.6400 88.6900 241.4000 ;
      RECT 87.5100 240.6400 87.8900 241.4000 ;
      RECT 86.7100 240.6400 87.0900 241.4000 ;
      RECT 85.9100 240.6400 86.2900 241.4000 ;
      RECT 85.1100 240.6400 85.4900 241.4000 ;
      RECT 84.3100 240.6400 84.6900 241.4000 ;
      RECT 83.5100 240.6400 83.8900 241.4000 ;
      RECT 82.7100 240.6400 83.0900 241.4000 ;
      RECT 81.9100 240.6400 82.2900 241.4000 ;
      RECT 81.1100 240.6400 81.4900 241.4000 ;
      RECT 80.3100 240.6400 80.6900 241.4000 ;
      RECT 79.5100 240.6400 79.8900 241.4000 ;
      RECT 78.7100 240.6400 79.0900 241.4000 ;
      RECT 77.9100 240.6400 78.2900 241.4000 ;
      RECT 77.1100 240.6400 77.4900 241.4000 ;
      RECT 76.3100 240.6400 76.6900 241.4000 ;
      RECT 75.5100 240.6400 75.8900 241.4000 ;
      RECT 74.7100 240.6400 75.0900 241.4000 ;
      RECT 73.9100 240.6400 74.2900 241.4000 ;
      RECT 73.1100 240.6400 73.4900 241.4000 ;
      RECT 72.3100 240.6400 72.6900 241.4000 ;
      RECT 71.5100 240.6400 71.8900 241.4000 ;
      RECT 70.7100 240.6400 71.0900 241.4000 ;
      RECT 69.9100 240.6400 70.2900 241.4000 ;
      RECT 69.1100 240.6400 69.4900 241.4000 ;
      RECT 68.3100 240.6400 68.6900 241.4000 ;
      RECT 67.5100 240.6400 67.8900 241.4000 ;
      RECT 66.7100 240.6400 67.0900 241.4000 ;
      RECT 65.9100 240.6400 66.2900 241.4000 ;
      RECT 65.1100 240.6400 65.4900 241.4000 ;
      RECT 64.3100 240.6400 64.6900 241.4000 ;
      RECT 63.5100 240.6400 63.8900 241.4000 ;
      RECT 62.7100 240.6400 63.0900 241.4000 ;
      RECT 61.9100 240.6400 62.2900 241.4000 ;
      RECT 61.1100 240.6400 61.4900 241.4000 ;
      RECT 60.3100 240.6400 60.6900 241.4000 ;
      RECT 59.5100 240.6400 59.8900 241.4000 ;
      RECT 58.7100 240.6400 59.0900 241.4000 ;
      RECT 57.9100 240.6400 58.2900 241.4000 ;
      RECT 0.0000 240.6400 57.4900 241.4000 ;
      RECT 0.0000 123.1500 243.0000 240.6400 ;
      RECT 0.7000 122.8500 243.0000 123.1500 ;
      RECT 0.0000 122.3500 243.0000 122.8500 ;
      RECT 0.7000 122.0500 243.0000 122.3500 ;
      RECT 0.0000 121.5500 243.0000 122.0500 ;
      RECT 0.7000 121.2500 243.0000 121.5500 ;
      RECT 0.0000 120.7500 243.0000 121.2500 ;
      RECT 0.7000 120.4500 243.0000 120.7500 ;
      RECT 0.0000 119.9500 243.0000 120.4500 ;
      RECT 0.7000 119.6500 243.0000 119.9500 ;
      RECT 0.0000 119.1500 243.0000 119.6500 ;
      RECT 0.7000 118.8500 243.0000 119.1500 ;
      RECT 0.0000 118.3500 243.0000 118.8500 ;
      RECT 0.7000 118.0500 243.0000 118.3500 ;
      RECT 0.0000 0.7600 243.0000 118.0500 ;
      RECT 185.1100 0.0000 243.0000 0.7600 ;
      RECT 184.3100 0.0000 184.6900 0.7600 ;
      RECT 183.5100 0.0000 183.8900 0.7600 ;
      RECT 182.7100 0.0000 183.0900 0.7600 ;
      RECT 181.9100 0.0000 182.2900 0.7600 ;
      RECT 181.1100 0.0000 181.4900 0.7600 ;
      RECT 180.3100 0.0000 180.6900 0.7600 ;
      RECT 179.5100 0.0000 179.8900 0.7600 ;
      RECT 178.7100 0.0000 179.0900 0.7600 ;
      RECT 177.9100 0.0000 178.2900 0.7600 ;
      RECT 177.1100 0.0000 177.4900 0.7600 ;
      RECT 176.3100 0.0000 176.6900 0.7600 ;
      RECT 175.5100 0.0000 175.8900 0.7600 ;
      RECT 174.7100 0.0000 175.0900 0.7600 ;
      RECT 173.9100 0.0000 174.2900 0.7600 ;
      RECT 173.1100 0.0000 173.4900 0.7600 ;
      RECT 172.3100 0.0000 172.6900 0.7600 ;
      RECT 171.5100 0.0000 171.8900 0.7600 ;
      RECT 170.7100 0.0000 171.0900 0.7600 ;
      RECT 169.9100 0.0000 170.2900 0.7600 ;
      RECT 169.1100 0.0000 169.4900 0.7600 ;
      RECT 168.3100 0.0000 168.6900 0.7600 ;
      RECT 167.5100 0.0000 167.8900 0.7600 ;
      RECT 166.7100 0.0000 167.0900 0.7600 ;
      RECT 165.9100 0.0000 166.2900 0.7600 ;
      RECT 165.1100 0.0000 165.4900 0.7600 ;
      RECT 164.3100 0.0000 164.6900 0.7600 ;
      RECT 163.5100 0.0000 163.8900 0.7600 ;
      RECT 162.7100 0.0000 163.0900 0.7600 ;
      RECT 161.9100 0.0000 162.2900 0.7600 ;
      RECT 161.1100 0.0000 161.4900 0.7600 ;
      RECT 160.3100 0.0000 160.6900 0.7600 ;
      RECT 159.5100 0.0000 159.8900 0.7600 ;
      RECT 158.7100 0.0000 159.0900 0.7600 ;
      RECT 157.9100 0.0000 158.2900 0.7600 ;
      RECT 157.1100 0.0000 157.4900 0.7600 ;
      RECT 156.3100 0.0000 156.6900 0.7600 ;
      RECT 155.5100 0.0000 155.8900 0.7600 ;
      RECT 154.7100 0.0000 155.0900 0.7600 ;
      RECT 153.9100 0.0000 154.2900 0.7600 ;
      RECT 153.1100 0.0000 153.4900 0.7600 ;
      RECT 152.3100 0.0000 152.6900 0.7600 ;
      RECT 151.5100 0.0000 151.8900 0.7600 ;
      RECT 150.7100 0.0000 151.0900 0.7600 ;
      RECT 149.9100 0.0000 150.2900 0.7600 ;
      RECT 149.1100 0.0000 149.4900 0.7600 ;
      RECT 148.3100 0.0000 148.6900 0.7600 ;
      RECT 147.5100 0.0000 147.8900 0.7600 ;
      RECT 146.7100 0.0000 147.0900 0.7600 ;
      RECT 145.9100 0.0000 146.2900 0.7600 ;
      RECT 145.1100 0.0000 145.4900 0.7600 ;
      RECT 144.3100 0.0000 144.6900 0.7600 ;
      RECT 143.5100 0.0000 143.8900 0.7600 ;
      RECT 142.7100 0.0000 143.0900 0.7600 ;
      RECT 141.9100 0.0000 142.2900 0.7600 ;
      RECT 141.1100 0.0000 141.4900 0.7600 ;
      RECT 140.3100 0.0000 140.6900 0.7600 ;
      RECT 139.5100 0.0000 139.8900 0.7600 ;
      RECT 138.7100 0.0000 139.0900 0.7600 ;
      RECT 137.9100 0.0000 138.2900 0.7600 ;
      RECT 137.1100 0.0000 137.4900 0.7600 ;
      RECT 136.3100 0.0000 136.6900 0.7600 ;
      RECT 135.5100 0.0000 135.8900 0.7600 ;
      RECT 134.7100 0.0000 135.0900 0.7600 ;
      RECT 133.9100 0.0000 134.2900 0.7600 ;
      RECT 133.1100 0.0000 133.4900 0.7600 ;
      RECT 132.3100 0.0000 132.6900 0.7600 ;
      RECT 131.5100 0.0000 131.8900 0.7600 ;
      RECT 130.7100 0.0000 131.0900 0.7600 ;
      RECT 129.9100 0.0000 130.2900 0.7600 ;
      RECT 129.1100 0.0000 129.4900 0.7600 ;
      RECT 128.3100 0.0000 128.6900 0.7600 ;
      RECT 127.5100 0.0000 127.8900 0.7600 ;
      RECT 126.7100 0.0000 127.0900 0.7600 ;
      RECT 125.9100 0.0000 126.2900 0.7600 ;
      RECT 125.1100 0.0000 125.4900 0.7600 ;
      RECT 124.3100 0.0000 124.6900 0.7600 ;
      RECT 123.5100 0.0000 123.8900 0.7600 ;
      RECT 122.7100 0.0000 123.0900 0.7600 ;
      RECT 121.9100 0.0000 122.2900 0.7600 ;
      RECT 121.1100 0.0000 121.4900 0.7600 ;
      RECT 120.3100 0.0000 120.6900 0.7600 ;
      RECT 119.5100 0.0000 119.8900 0.7600 ;
      RECT 118.7100 0.0000 119.0900 0.7600 ;
      RECT 117.9100 0.0000 118.2900 0.7600 ;
      RECT 117.1100 0.0000 117.4900 0.7600 ;
      RECT 116.3100 0.0000 116.6900 0.7600 ;
      RECT 115.5100 0.0000 115.8900 0.7600 ;
      RECT 114.7100 0.0000 115.0900 0.7600 ;
      RECT 113.9100 0.0000 114.2900 0.7600 ;
      RECT 113.1100 0.0000 113.4900 0.7600 ;
      RECT 112.3100 0.0000 112.6900 0.7600 ;
      RECT 111.5100 0.0000 111.8900 0.7600 ;
      RECT 110.7100 0.0000 111.0900 0.7600 ;
      RECT 109.9100 0.0000 110.2900 0.7600 ;
      RECT 109.1100 0.0000 109.4900 0.7600 ;
      RECT 108.3100 0.0000 108.6900 0.7600 ;
      RECT 107.5100 0.0000 107.8900 0.7600 ;
      RECT 106.7100 0.0000 107.0900 0.7600 ;
      RECT 105.9100 0.0000 106.2900 0.7600 ;
      RECT 105.1100 0.0000 105.4900 0.7600 ;
      RECT 104.3100 0.0000 104.6900 0.7600 ;
      RECT 103.5100 0.0000 103.8900 0.7600 ;
      RECT 102.7100 0.0000 103.0900 0.7600 ;
      RECT 101.9100 0.0000 102.2900 0.7600 ;
      RECT 101.1100 0.0000 101.4900 0.7600 ;
      RECT 100.3100 0.0000 100.6900 0.7600 ;
      RECT 99.5100 0.0000 99.8900 0.7600 ;
      RECT 98.7100 0.0000 99.0900 0.7600 ;
      RECT 97.9100 0.0000 98.2900 0.7600 ;
      RECT 97.1100 0.0000 97.4900 0.7600 ;
      RECT 96.3100 0.0000 96.6900 0.7600 ;
      RECT 95.5100 0.0000 95.8900 0.7600 ;
      RECT 94.7100 0.0000 95.0900 0.7600 ;
      RECT 93.9100 0.0000 94.2900 0.7600 ;
      RECT 93.1100 0.0000 93.4900 0.7600 ;
      RECT 92.3100 0.0000 92.6900 0.7600 ;
      RECT 91.5100 0.0000 91.8900 0.7600 ;
      RECT 90.7100 0.0000 91.0900 0.7600 ;
      RECT 89.9100 0.0000 90.2900 0.7600 ;
      RECT 89.1100 0.0000 89.4900 0.7600 ;
      RECT 88.3100 0.0000 88.6900 0.7600 ;
      RECT 87.5100 0.0000 87.8900 0.7600 ;
      RECT 86.7100 0.0000 87.0900 0.7600 ;
      RECT 85.9100 0.0000 86.2900 0.7600 ;
      RECT 85.1100 0.0000 85.4900 0.7600 ;
      RECT 84.3100 0.0000 84.6900 0.7600 ;
      RECT 83.5100 0.0000 83.8900 0.7600 ;
      RECT 82.7100 0.0000 83.0900 0.7600 ;
      RECT 81.9100 0.0000 82.2900 0.7600 ;
      RECT 81.1100 0.0000 81.4900 0.7600 ;
      RECT 80.3100 0.0000 80.6900 0.7600 ;
      RECT 79.5100 0.0000 79.8900 0.7600 ;
      RECT 78.7100 0.0000 79.0900 0.7600 ;
      RECT 77.9100 0.0000 78.2900 0.7600 ;
      RECT 77.1100 0.0000 77.4900 0.7600 ;
      RECT 76.3100 0.0000 76.6900 0.7600 ;
      RECT 75.5100 0.0000 75.8900 0.7600 ;
      RECT 74.7100 0.0000 75.0900 0.7600 ;
      RECT 73.9100 0.0000 74.2900 0.7600 ;
      RECT 73.1100 0.0000 73.4900 0.7600 ;
      RECT 72.3100 0.0000 72.6900 0.7600 ;
      RECT 71.5100 0.0000 71.8900 0.7600 ;
      RECT 70.7100 0.0000 71.0900 0.7600 ;
      RECT 69.9100 0.0000 70.2900 0.7600 ;
      RECT 69.1100 0.0000 69.4900 0.7600 ;
      RECT 68.3100 0.0000 68.6900 0.7600 ;
      RECT 67.5100 0.0000 67.8900 0.7600 ;
      RECT 66.7100 0.0000 67.0900 0.7600 ;
      RECT 65.9100 0.0000 66.2900 0.7600 ;
      RECT 65.1100 0.0000 65.4900 0.7600 ;
      RECT 64.3100 0.0000 64.6900 0.7600 ;
      RECT 63.5100 0.0000 63.8900 0.7600 ;
      RECT 62.7100 0.0000 63.0900 0.7600 ;
      RECT 61.9100 0.0000 62.2900 0.7600 ;
      RECT 61.1100 0.0000 61.4900 0.7600 ;
      RECT 60.3100 0.0000 60.6900 0.7600 ;
      RECT 59.5100 0.0000 59.8900 0.7600 ;
      RECT 58.7100 0.0000 59.0900 0.7600 ;
      RECT 57.9100 0.0000 58.2900 0.7600 ;
      RECT 0.0000 0.0000 57.4900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 240.7250 243.0000 241.4000 ;
      RECT 240.1600 240.5600 243.0000 240.7250 ;
      RECT 2.1600 240.5600 238.8400 240.7250 ;
      RECT 240.1600 0.8400 240.8400 240.5600 ;
      RECT 4.1600 0.8400 238.8400 240.5600 ;
      RECT 2.1600 0.8400 2.8400 240.5600 ;
      RECT 0.0000 0.8400 0.8400 240.7250 ;
      RECT 242.1600 0.6750 243.0000 240.5600 ;
      RECT 4.1600 0.6750 240.8400 0.8400 ;
      RECT 0.0000 0.6750 2.8400 0.8400 ;
      RECT 0.0000 0.0000 243.0000 0.6750 ;
  END
END sram_160b_w16

END LIBRARY
