##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sun Mar  9 21:32:38 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 479.0000 BY 477.2000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 192.7500 0.6000 192.8500 ;
    END
  END clk
  PIN sum_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.2500 0.0000 239.3500 0.6000 ;
    END
  END sum_out[159]
  PIN sum_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 238.2500 0.0000 238.3500 0.6000 ;
    END
  END sum_out[158]
  PIN sum_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 237.2500 0.0000 237.3500 0.6000 ;
    END
  END sum_out[157]
  PIN sum_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.2500 0.0000 236.3500 0.6000 ;
    END
  END sum_out[156]
  PIN sum_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 235.2500 0.0000 235.3500 0.6000 ;
    END
  END sum_out[155]
  PIN sum_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 234.2500 0.0000 234.3500 0.6000 ;
    END
  END sum_out[154]
  PIN sum_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.2500 0.0000 233.3500 0.6000 ;
    END
  END sum_out[153]
  PIN sum_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 232.2500 0.0000 232.3500 0.6000 ;
    END
  END sum_out[152]
  PIN sum_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.2500 0.0000 231.3500 0.6000 ;
    END
  END sum_out[151]
  PIN sum_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 230.2500 0.0000 230.3500 0.6000 ;
    END
  END sum_out[150]
  PIN sum_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 229.2500 0.0000 229.3500 0.6000 ;
    END
  END sum_out[149]
  PIN sum_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.2500 0.0000 228.3500 0.6000 ;
    END
  END sum_out[148]
  PIN sum_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 227.2500 0.0000 227.3500 0.6000 ;
    END
  END sum_out[147]
  PIN sum_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.2500 0.0000 226.3500 0.6000 ;
    END
  END sum_out[146]
  PIN sum_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.2500 0.0000 225.3500 0.6000 ;
    END
  END sum_out[145]
  PIN sum_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 224.2500 0.0000 224.3500 0.6000 ;
    END
  END sum_out[144]
  PIN sum_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.2500 0.0000 223.3500 0.6000 ;
    END
  END sum_out[143]
  PIN sum_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 222.2500 0.0000 222.3500 0.6000 ;
    END
  END sum_out[142]
  PIN sum_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.2500 0.0000 221.3500 0.6000 ;
    END
  END sum_out[141]
  PIN sum_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.2500 0.0000 220.3500 0.6000 ;
    END
  END sum_out[140]
  PIN sum_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 219.2500 0.0000 219.3500 0.6000 ;
    END
  END sum_out[139]
  PIN sum_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.2500 0.0000 218.3500 0.6000 ;
    END
  END sum_out[138]
  PIN sum_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.2500 0.0000 217.3500 0.6000 ;
    END
  END sum_out[137]
  PIN sum_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 216.2500 0.0000 216.3500 0.6000 ;
    END
  END sum_out[136]
  PIN sum_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.2500 0.0000 215.3500 0.6000 ;
    END
  END sum_out[135]
  PIN sum_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 214.2500 0.0000 214.3500 0.6000 ;
    END
  END sum_out[134]
  PIN sum_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.2500 0.0000 213.3500 0.6000 ;
    END
  END sum_out[133]
  PIN sum_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.2500 0.0000 212.3500 0.6000 ;
    END
  END sum_out[132]
  PIN sum_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 211.2500 0.0000 211.3500 0.6000 ;
    END
  END sum_out[131]
  PIN sum_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.2500 0.0000 210.3500 0.6000 ;
    END
  END sum_out[130]
  PIN sum_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.2500 0.0000 209.3500 0.6000 ;
    END
  END sum_out[129]
  PIN sum_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 208.2500 0.0000 208.3500 0.6000 ;
    END
  END sum_out[128]
  PIN sum_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.2500 0.0000 207.3500 0.6000 ;
    END
  END sum_out[127]
  PIN sum_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 206.2500 0.0000 206.3500 0.6000 ;
    END
  END sum_out[126]
  PIN sum_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.2500 0.0000 205.3500 0.6000 ;
    END
  END sum_out[125]
  PIN sum_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.2500 0.0000 204.3500 0.6000 ;
    END
  END sum_out[124]
  PIN sum_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 203.2500 0.0000 203.3500 0.6000 ;
    END
  END sum_out[123]
  PIN sum_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.2500 0.0000 202.3500 0.6000 ;
    END
  END sum_out[122]
  PIN sum_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.2500 0.0000 201.3500 0.6000 ;
    END
  END sum_out[121]
  PIN sum_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 200.2500 0.0000 200.3500 0.6000 ;
    END
  END sum_out[120]
  PIN sum_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.2500 0.0000 199.3500 0.6000 ;
    END
  END sum_out[119]
  PIN sum_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 198.2500 0.0000 198.3500 0.6000 ;
    END
  END sum_out[118]
  PIN sum_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.2500 0.0000 197.3500 0.6000 ;
    END
  END sum_out[117]
  PIN sum_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.2500 0.0000 196.3500 0.6000 ;
    END
  END sum_out[116]
  PIN sum_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 195.2500 0.0000 195.3500 0.6000 ;
    END
  END sum_out[115]
  PIN sum_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.2500 0.0000 194.3500 0.6000 ;
    END
  END sum_out[114]
  PIN sum_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.2500 0.0000 193.3500 0.6000 ;
    END
  END sum_out[113]
  PIN sum_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 192.2500 0.0000 192.3500 0.6000 ;
    END
  END sum_out[112]
  PIN sum_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.2500 0.0000 191.3500 0.6000 ;
    END
  END sum_out[111]
  PIN sum_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 190.2500 0.0000 190.3500 0.6000 ;
    END
  END sum_out[110]
  PIN sum_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.2500 0.0000 189.3500 0.6000 ;
    END
  END sum_out[109]
  PIN sum_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.2500 0.0000 188.3500 0.6000 ;
    END
  END sum_out[108]
  PIN sum_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 187.2500 0.0000 187.3500 0.6000 ;
    END
  END sum_out[107]
  PIN sum_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.2500 0.0000 186.3500 0.6000 ;
    END
  END sum_out[106]
  PIN sum_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.2500 0.0000 185.3500 0.6000 ;
    END
  END sum_out[105]
  PIN sum_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.2500 0.0000 184.3500 0.6000 ;
    END
  END sum_out[104]
  PIN sum_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.2500 0.0000 183.3500 0.6000 ;
    END
  END sum_out[103]
  PIN sum_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.2500 0.0000 182.3500 0.6000 ;
    END
  END sum_out[102]
  PIN sum_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.2500 0.0000 181.3500 0.6000 ;
    END
  END sum_out[101]
  PIN sum_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.2500 0.0000 180.3500 0.6000 ;
    END
  END sum_out[100]
  PIN sum_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.2500 0.0000 179.3500 0.6000 ;
    END
  END sum_out[99]
  PIN sum_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.2500 0.0000 178.3500 0.6000 ;
    END
  END sum_out[98]
  PIN sum_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.2500 0.0000 177.3500 0.6000 ;
    END
  END sum_out[97]
  PIN sum_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.2500 0.0000 176.3500 0.6000 ;
    END
  END sum_out[96]
  PIN sum_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.2500 0.0000 175.3500 0.6000 ;
    END
  END sum_out[95]
  PIN sum_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.2500 0.0000 174.3500 0.6000 ;
    END
  END sum_out[94]
  PIN sum_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.2500 0.0000 173.3500 0.6000 ;
    END
  END sum_out[93]
  PIN sum_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.2500 0.0000 172.3500 0.6000 ;
    END
  END sum_out[92]
  PIN sum_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.2500 0.0000 171.3500 0.6000 ;
    END
  END sum_out[91]
  PIN sum_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.2500 0.0000 170.3500 0.6000 ;
    END
  END sum_out[90]
  PIN sum_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.2500 0.0000 169.3500 0.6000 ;
    END
  END sum_out[89]
  PIN sum_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.2500 0.0000 168.3500 0.6000 ;
    END
  END sum_out[88]
  PIN sum_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.2500 0.0000 167.3500 0.6000 ;
    END
  END sum_out[87]
  PIN sum_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.2500 0.0000 166.3500 0.6000 ;
    END
  END sum_out[86]
  PIN sum_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.2500 0.0000 165.3500 0.6000 ;
    END
  END sum_out[85]
  PIN sum_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.2500 0.0000 164.3500 0.6000 ;
    END
  END sum_out[84]
  PIN sum_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.2500 0.0000 163.3500 0.6000 ;
    END
  END sum_out[83]
  PIN sum_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.2500 0.0000 162.3500 0.6000 ;
    END
  END sum_out[82]
  PIN sum_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.2500 0.0000 161.3500 0.6000 ;
    END
  END sum_out[81]
  PIN sum_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.2500 0.0000 160.3500 0.6000 ;
    END
  END sum_out[80]
  PIN sum_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.2500 0.0000 159.3500 0.6000 ;
    END
  END sum_out[79]
  PIN sum_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.2500 0.0000 158.3500 0.6000 ;
    END
  END sum_out[78]
  PIN sum_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.2500 0.0000 157.3500 0.6000 ;
    END
  END sum_out[77]
  PIN sum_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.2500 0.0000 156.3500 0.6000 ;
    END
  END sum_out[76]
  PIN sum_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.2500 0.0000 155.3500 0.6000 ;
    END
  END sum_out[75]
  PIN sum_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.2500 0.0000 154.3500 0.6000 ;
    END
  END sum_out[74]
  PIN sum_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.2500 0.0000 153.3500 0.6000 ;
    END
  END sum_out[73]
  PIN sum_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.2500 0.0000 152.3500 0.6000 ;
    END
  END sum_out[72]
  PIN sum_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.2500 0.0000 151.3500 0.6000 ;
    END
  END sum_out[71]
  PIN sum_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.2500 0.0000 150.3500 0.6000 ;
    END
  END sum_out[70]
  PIN sum_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.2500 0.0000 149.3500 0.6000 ;
    END
  END sum_out[69]
  PIN sum_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.2500 0.0000 148.3500 0.6000 ;
    END
  END sum_out[68]
  PIN sum_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.2500 0.0000 147.3500 0.6000 ;
    END
  END sum_out[67]
  PIN sum_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.2500 0.0000 146.3500 0.6000 ;
    END
  END sum_out[66]
  PIN sum_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.2500 0.0000 145.3500 0.6000 ;
    END
  END sum_out[65]
  PIN sum_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.2500 0.0000 144.3500 0.6000 ;
    END
  END sum_out[64]
  PIN sum_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.2500 0.0000 143.3500 0.6000 ;
    END
  END sum_out[63]
  PIN sum_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 142.2500 0.0000 142.3500 0.6000 ;
    END
  END sum_out[62]
  PIN sum_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.2500 0.0000 141.3500 0.6000 ;
    END
  END sum_out[61]
  PIN sum_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.2500 0.0000 140.3500 0.6000 ;
    END
  END sum_out[60]
  PIN sum_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 139.2500 0.0000 139.3500 0.6000 ;
    END
  END sum_out[59]
  PIN sum_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.2500 0.0000 138.3500 0.6000 ;
    END
  END sum_out[58]
  PIN sum_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.2500 0.0000 137.3500 0.6000 ;
    END
  END sum_out[57]
  PIN sum_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.2500 0.0000 136.3500 0.6000 ;
    END
  END sum_out[56]
  PIN sum_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.2500 0.0000 135.3500 0.6000 ;
    END
  END sum_out[55]
  PIN sum_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.2500 0.0000 134.3500 0.6000 ;
    END
  END sum_out[54]
  PIN sum_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.2500 0.0000 133.3500 0.6000 ;
    END
  END sum_out[53]
  PIN sum_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.2500 0.0000 132.3500 0.6000 ;
    END
  END sum_out[52]
  PIN sum_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.2500 0.0000 131.3500 0.6000 ;
    END
  END sum_out[51]
  PIN sum_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.2500 0.0000 130.3500 0.6000 ;
    END
  END sum_out[50]
  PIN sum_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.2500 0.0000 129.3500 0.6000 ;
    END
  END sum_out[49]
  PIN sum_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.2500 0.0000 128.3500 0.6000 ;
    END
  END sum_out[48]
  PIN sum_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.2500 0.0000 127.3500 0.6000 ;
    END
  END sum_out[47]
  PIN sum_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 126.2500 0.0000 126.3500 0.6000 ;
    END
  END sum_out[46]
  PIN sum_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.2500 0.0000 125.3500 0.6000 ;
    END
  END sum_out[45]
  PIN sum_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.2500 0.0000 124.3500 0.6000 ;
    END
  END sum_out[44]
  PIN sum_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.2500 0.0000 123.3500 0.6000 ;
    END
  END sum_out[43]
  PIN sum_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.2500 0.0000 122.3500 0.6000 ;
    END
  END sum_out[42]
  PIN sum_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.2500 0.0000 121.3500 0.6000 ;
    END
  END sum_out[41]
  PIN sum_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.2500 0.0000 120.3500 0.6000 ;
    END
  END sum_out[40]
  PIN sum_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.2500 0.0000 119.3500 0.6000 ;
    END
  END sum_out[39]
  PIN sum_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 118.2500 0.0000 118.3500 0.6000 ;
    END
  END sum_out[38]
  PIN sum_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.2500 0.0000 117.3500 0.6000 ;
    END
  END sum_out[37]
  PIN sum_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.2500 0.0000 116.3500 0.6000 ;
    END
  END sum_out[36]
  PIN sum_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.2500 0.0000 115.3500 0.6000 ;
    END
  END sum_out[35]
  PIN sum_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.2500 0.0000 114.3500 0.6000 ;
    END
  END sum_out[34]
  PIN sum_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.2500 0.0000 113.3500 0.6000 ;
    END
  END sum_out[33]
  PIN sum_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.2500 0.0000 112.3500 0.6000 ;
    END
  END sum_out[32]
  PIN sum_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.2500 0.0000 111.3500 0.6000 ;
    END
  END sum_out[31]
  PIN sum_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 110.2500 0.0000 110.3500 0.6000 ;
    END
  END sum_out[30]
  PIN sum_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.2500 0.0000 109.3500 0.6000 ;
    END
  END sum_out[29]
  PIN sum_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.2500 0.0000 108.3500 0.6000 ;
    END
  END sum_out[28]
  PIN sum_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 107.2500 0.0000 107.3500 0.6000 ;
    END
  END sum_out[27]
  PIN sum_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.2500 0.0000 106.3500 0.6000 ;
    END
  END sum_out[26]
  PIN sum_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.2500 0.0000 105.3500 0.6000 ;
    END
  END sum_out[25]
  PIN sum_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.2500 0.0000 104.3500 0.6000 ;
    END
  END sum_out[24]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.2500 0.0000 103.3500 0.6000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 102.2500 0.0000 102.3500 0.6000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.2500 0.0000 101.3500 0.6000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.2500 0.0000 100.3500 0.6000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 99.2500 0.0000 99.3500 0.6000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.2500 0.0000 98.3500 0.6000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.2500 0.0000 97.3500 0.6000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.2500 0.0000 96.3500 0.6000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.2500 0.0000 95.3500 0.6000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 94.2500 0.0000 94.3500 0.6000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.2500 0.0000 93.3500 0.6000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.2500 0.0000 92.3500 0.6000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.2500 0.0000 91.3500 0.6000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.2500 0.0000 90.3500 0.6000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.2500 0.0000 89.3500 0.6000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.2500 0.0000 88.3500 0.6000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.2500 0.0000 87.3500 0.6000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.2500 0.0000 86.3500 0.6000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.2500 0.0000 85.3500 0.6000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.2500 0.0000 84.3500 0.6000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 83.2500 0.0000 83.3500 0.6000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.2500 0.0000 82.3500 0.6000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.2500 0.0000 81.3500 0.6000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.2500 0.0000 80.3500 0.6000 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 320.7500 0.6000 320.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 318.7500 0.6000 318.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 316.7500 0.6000 316.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 314.7500 0.6000 314.8500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 312.7500 0.6000 312.8500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 310.7500 0.6000 310.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 308.7500 0.6000 308.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 306.7500 0.6000 306.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 304.7500 0.6000 304.8500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 302.7500 0.6000 302.8500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 300.7500 0.6000 300.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 298.7500 0.6000 298.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 296.7500 0.6000 296.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 294.7500 0.6000 294.8500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 292.7500 0.6000 292.8500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 290.7500 0.6000 290.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 288.7500 0.6000 288.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 286.7500 0.6000 286.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 284.7500 0.6000 284.8500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 282.7500 0.6000 282.8500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 280.7500 0.6000 280.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 278.7500 0.6000 278.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 276.7500 0.6000 276.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 274.7500 0.6000 274.8500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 272.7500 0.6000 272.8500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 270.7500 0.6000 270.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 268.7500 0.6000 268.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 266.7500 0.6000 266.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 264.7500 0.6000 264.8500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 262.7500 0.6000 262.8500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 260.7500 0.6000 260.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 258.7500 0.6000 258.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 256.7500 0.6000 256.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 254.7500 0.6000 254.8500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 252.7500 0.6000 252.8500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 250.7500 0.6000 250.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 248.7500 0.6000 248.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 246.7500 0.6000 246.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 244.7500 0.6000 244.8500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 242.7500 0.6000 242.8500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 240.7500 0.6000 240.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 238.7500 0.6000 238.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 236.7500 0.6000 236.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 234.7500 0.6000 234.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 232.7500 0.6000 232.8500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 230.7500 0.6000 230.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 228.7500 0.6000 228.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 226.7500 0.6000 226.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 224.7500 0.6000 224.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 222.7500 0.6000 222.8500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 220.7500 0.6000 220.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 218.7500 0.6000 218.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 216.7500 0.6000 216.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 214.7500 0.6000 214.8500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 212.7500 0.6000 212.8500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.7500 0.6000 210.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 208.7500 0.6000 208.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 206.7500 0.6000 206.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 204.7500 0.6000 204.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 202.7500 0.6000 202.8500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 200.7500 0.6000 200.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.7500 0.6000 198.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 196.7500 0.6000 196.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 194.7500 0.6000 194.8500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 399.2500 0.0000 399.3500 0.6000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 398.2500 0.0000 398.3500 0.6000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 397.2500 0.0000 397.3500 0.6000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 396.2500 0.0000 396.3500 0.6000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 395.2500 0.0000 395.3500 0.6000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 394.2500 0.0000 394.3500 0.6000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 393.2500 0.0000 393.3500 0.6000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 392.2500 0.0000 392.3500 0.6000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 391.2500 0.0000 391.3500 0.6000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 390.2500 0.0000 390.3500 0.6000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.2500 0.0000 389.3500 0.6000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 388.2500 0.0000 388.3500 0.6000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 387.2500 0.0000 387.3500 0.6000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.2500 0.0000 386.3500 0.6000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 385.2500 0.0000 385.3500 0.6000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 384.2500 0.0000 384.3500 0.6000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.2500 0.0000 383.3500 0.6000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.2500 0.0000 382.3500 0.6000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 381.2500 0.0000 381.3500 0.6000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.2500 0.0000 380.3500 0.6000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 379.2500 0.0000 379.3500 0.6000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.2500 0.0000 378.3500 0.6000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.2500 0.0000 377.3500 0.6000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 376.2500 0.0000 376.3500 0.6000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.2500 0.0000 375.3500 0.6000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 374.2500 0.0000 374.3500 0.6000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 373.2500 0.0000 373.3500 0.6000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.2500 0.0000 372.3500 0.6000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 371.2500 0.0000 371.3500 0.6000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.2500 0.0000 370.3500 0.6000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 369.2500 0.0000 369.3500 0.6000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 368.2500 0.0000 368.3500 0.6000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.2500 0.0000 367.3500 0.6000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 366.2500 0.0000 366.3500 0.6000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.2500 0.0000 365.3500 0.6000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 364.2500 0.0000 364.3500 0.6000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.2500 0.0000 363.3500 0.6000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.2500 0.0000 362.3500 0.6000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 361.2500 0.0000 361.3500 0.6000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 360.2500 0.0000 360.3500 0.6000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.2500 0.0000 359.3500 0.6000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 358.2500 0.0000 358.3500 0.6000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.2500 0.0000 357.3500 0.6000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 356.2500 0.0000 356.3500 0.6000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 355.2500 0.0000 355.3500 0.6000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.2500 0.0000 354.3500 0.6000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.2500 0.0000 353.3500 0.6000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 352.2500 0.0000 352.3500 0.6000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.2500 0.0000 351.3500 0.6000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 350.2500 0.0000 350.3500 0.6000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 349.2500 0.0000 349.3500 0.6000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.2500 0.0000 348.3500 0.6000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 347.2500 0.0000 347.3500 0.6000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.2500 0.0000 346.3500 0.6000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.2500 0.0000 345.3500 0.6000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 344.2500 0.0000 344.3500 0.6000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.2500 0.0000 343.3500 0.6000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.2500 0.0000 342.3500 0.6000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.2500 0.0000 341.3500 0.6000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.2500 0.0000 340.3500 0.6000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.2500 0.0000 339.3500 0.6000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.2500 0.0000 338.3500 0.6000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.2500 0.0000 337.3500 0.6000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.2500 0.0000 336.3500 0.6000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.2500 0.0000 335.3500 0.6000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.2500 0.0000 334.3500 0.6000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.2500 0.0000 333.3500 0.6000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.2500 0.0000 332.3500 0.6000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.2500 0.0000 331.3500 0.6000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.2500 0.0000 330.3500 0.6000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.2500 0.0000 329.3500 0.6000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 328.2500 0.0000 328.3500 0.6000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.2500 0.0000 327.3500 0.6000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 326.2500 0.0000 326.3500 0.6000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.2500 0.0000 325.3500 0.6000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.2500 0.0000 324.3500 0.6000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.2500 0.0000 323.3500 0.6000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.2500 0.0000 322.3500 0.6000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.2500 0.0000 321.3500 0.6000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 320.2500 0.0000 320.3500 0.6000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.2500 0.0000 319.3500 0.6000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.2500 0.0000 318.3500 0.6000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.2500 0.0000 317.3500 0.6000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.2500 0.0000 316.3500 0.6000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.2500 0.0000 315.3500 0.6000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.2500 0.0000 314.3500 0.6000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.2500 0.0000 313.3500 0.6000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.2500 0.0000 312.3500 0.6000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.2500 0.0000 311.3500 0.6000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.2500 0.0000 310.3500 0.6000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.2500 0.0000 309.3500 0.6000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.2500 0.0000 308.3500 0.6000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.2500 0.0000 307.3500 0.6000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.2500 0.0000 306.3500 0.6000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.2500 0.0000 305.3500 0.6000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 304.2500 0.0000 304.3500 0.6000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.2500 0.0000 303.3500 0.6000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 302.2500 0.0000 302.3500 0.6000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.2500 0.0000 301.3500 0.6000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.2500 0.0000 300.3500 0.6000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.2500 0.0000 299.3500 0.6000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.2500 0.0000 298.3500 0.6000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.2500 0.0000 297.3500 0.6000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 296.2500 0.0000 296.3500 0.6000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.2500 0.0000 295.3500 0.6000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 294.2500 0.0000 294.3500 0.6000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.2500 0.0000 293.3500 0.6000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.2500 0.0000 292.3500 0.6000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.2500 0.0000 291.3500 0.6000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.2500 0.0000 290.3500 0.6000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.2500 0.0000 289.3500 0.6000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 288.2500 0.0000 288.3500 0.6000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.2500 0.0000 287.3500 0.6000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.2500 0.0000 286.3500 0.6000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 285.2500 0.0000 285.3500 0.6000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 284.2500 0.0000 284.3500 0.6000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.2500 0.0000 283.3500 0.6000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.2500 0.0000 282.3500 0.6000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.2500 0.0000 281.3500 0.6000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 280.2500 0.0000 280.3500 0.6000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.2500 0.0000 279.3500 0.6000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 278.2500 0.0000 278.3500 0.6000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.2500 0.0000 277.3500 0.6000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.2500 0.0000 276.3500 0.6000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 275.2500 0.0000 275.3500 0.6000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.2500 0.0000 274.3500 0.6000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 273.2500 0.0000 273.3500 0.6000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 272.2500 0.0000 272.3500 0.6000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.2500 0.0000 271.3500 0.6000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 270.2500 0.0000 270.3500 0.6000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 269.2500 0.0000 269.3500 0.6000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 268.2500 0.0000 268.3500 0.6000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 267.2500 0.0000 267.3500 0.6000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 266.2500 0.0000 266.3500 0.6000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 265.2500 0.0000 265.3500 0.6000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 264.2500 0.0000 264.3500 0.6000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 263.2500 0.0000 263.3500 0.6000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 262.2500 0.0000 262.3500 0.6000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 261.2500 0.0000 261.3500 0.6000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 260.2500 0.0000 260.3500 0.6000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 259.2500 0.0000 259.3500 0.6000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 258.2500 0.0000 258.3500 0.6000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 257.2500 0.0000 257.3500 0.6000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 256.2500 0.0000 256.3500 0.6000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.2500 0.0000 255.3500 0.6000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 254.2500 0.0000 254.3500 0.6000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 253.2500 0.0000 253.3500 0.6000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.2500 0.0000 252.3500 0.6000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 251.2500 0.0000 251.3500 0.6000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.2500 0.0000 250.3500 0.6000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 249.2500 0.0000 249.3500 0.6000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 248.2500 0.0000 248.3500 0.6000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.2500 0.0000 247.3500 0.6000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 246.2500 0.0000 246.3500 0.6000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.2500 0.0000 245.3500 0.6000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.2500 0.0000 244.3500 0.6000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 243.2500 0.0000 243.3500 0.6000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.2500 0.0000 242.3500 0.6000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 241.2500 0.0000 241.3500 0.6000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 240.2500 0.0000 240.3500 0.6000 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 190.7500 0.6000 190.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 188.7500 0.6000 188.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.7500 0.6000 186.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 184.7500 0.6000 184.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 182.7500 0.6000 182.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 180.7500 0.6000 180.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 178.7500 0.6000 178.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 176.7500 0.6000 176.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 174.7500 0.6000 174.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 172.7500 0.6000 172.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 170.7500 0.6000 170.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 168.7500 0.6000 168.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 166.7500 0.6000 166.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 164.7500 0.6000 164.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 162.7500 0.6000 162.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 160.7500 0.6000 160.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 158.7500 0.6000 158.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 156.7500 0.6000 156.8500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
    LAYER M3 ;
      RECT 0.0000 320.9500 479.0000 477.2000 ;
      RECT 0.7000 320.6500 479.0000 320.9500 ;
      RECT 0.0000 318.9500 479.0000 320.6500 ;
      RECT 0.7000 318.6500 479.0000 318.9500 ;
      RECT 0.0000 316.9500 479.0000 318.6500 ;
      RECT 0.7000 316.6500 479.0000 316.9500 ;
      RECT 0.0000 314.9500 479.0000 316.6500 ;
      RECT 0.7000 314.6500 479.0000 314.9500 ;
      RECT 0.0000 312.9500 479.0000 314.6500 ;
      RECT 0.7000 312.6500 479.0000 312.9500 ;
      RECT 0.0000 310.9500 479.0000 312.6500 ;
      RECT 0.7000 310.6500 479.0000 310.9500 ;
      RECT 0.0000 308.9500 479.0000 310.6500 ;
      RECT 0.7000 308.6500 479.0000 308.9500 ;
      RECT 0.0000 306.9500 479.0000 308.6500 ;
      RECT 0.7000 306.6500 479.0000 306.9500 ;
      RECT 0.0000 304.9500 479.0000 306.6500 ;
      RECT 0.7000 304.6500 479.0000 304.9500 ;
      RECT 0.0000 302.9500 479.0000 304.6500 ;
      RECT 0.7000 302.6500 479.0000 302.9500 ;
      RECT 0.0000 300.9500 479.0000 302.6500 ;
      RECT 0.7000 300.6500 479.0000 300.9500 ;
      RECT 0.0000 298.9500 479.0000 300.6500 ;
      RECT 0.7000 298.6500 479.0000 298.9500 ;
      RECT 0.0000 296.9500 479.0000 298.6500 ;
      RECT 0.7000 296.6500 479.0000 296.9500 ;
      RECT 0.0000 294.9500 479.0000 296.6500 ;
      RECT 0.7000 294.6500 479.0000 294.9500 ;
      RECT 0.0000 292.9500 479.0000 294.6500 ;
      RECT 0.7000 292.6500 479.0000 292.9500 ;
      RECT 0.0000 290.9500 479.0000 292.6500 ;
      RECT 0.7000 290.6500 479.0000 290.9500 ;
      RECT 0.0000 288.9500 479.0000 290.6500 ;
      RECT 0.7000 288.6500 479.0000 288.9500 ;
      RECT 0.0000 286.9500 479.0000 288.6500 ;
      RECT 0.7000 286.6500 479.0000 286.9500 ;
      RECT 0.0000 284.9500 479.0000 286.6500 ;
      RECT 0.7000 284.6500 479.0000 284.9500 ;
      RECT 0.0000 282.9500 479.0000 284.6500 ;
      RECT 0.7000 282.6500 479.0000 282.9500 ;
      RECT 0.0000 280.9500 479.0000 282.6500 ;
      RECT 0.7000 280.6500 479.0000 280.9500 ;
      RECT 0.0000 278.9500 479.0000 280.6500 ;
      RECT 0.7000 278.6500 479.0000 278.9500 ;
      RECT 0.0000 276.9500 479.0000 278.6500 ;
      RECT 0.7000 276.6500 479.0000 276.9500 ;
      RECT 0.0000 274.9500 479.0000 276.6500 ;
      RECT 0.7000 274.6500 479.0000 274.9500 ;
      RECT 0.0000 272.9500 479.0000 274.6500 ;
      RECT 0.7000 272.6500 479.0000 272.9500 ;
      RECT 0.0000 270.9500 479.0000 272.6500 ;
      RECT 0.7000 270.6500 479.0000 270.9500 ;
      RECT 0.0000 268.9500 479.0000 270.6500 ;
      RECT 0.7000 268.6500 479.0000 268.9500 ;
      RECT 0.0000 266.9500 479.0000 268.6500 ;
      RECT 0.7000 266.6500 479.0000 266.9500 ;
      RECT 0.0000 264.9500 479.0000 266.6500 ;
      RECT 0.7000 264.6500 479.0000 264.9500 ;
      RECT 0.0000 262.9500 479.0000 264.6500 ;
      RECT 0.7000 262.6500 479.0000 262.9500 ;
      RECT 0.0000 260.9500 479.0000 262.6500 ;
      RECT 0.7000 260.6500 479.0000 260.9500 ;
      RECT 0.0000 258.9500 479.0000 260.6500 ;
      RECT 0.7000 258.6500 479.0000 258.9500 ;
      RECT 0.0000 256.9500 479.0000 258.6500 ;
      RECT 0.7000 256.6500 479.0000 256.9500 ;
      RECT 0.0000 254.9500 479.0000 256.6500 ;
      RECT 0.7000 254.6500 479.0000 254.9500 ;
      RECT 0.0000 252.9500 479.0000 254.6500 ;
      RECT 0.7000 252.6500 479.0000 252.9500 ;
      RECT 0.0000 250.9500 479.0000 252.6500 ;
      RECT 0.7000 250.6500 479.0000 250.9500 ;
      RECT 0.0000 248.9500 479.0000 250.6500 ;
      RECT 0.7000 248.6500 479.0000 248.9500 ;
      RECT 0.0000 246.9500 479.0000 248.6500 ;
      RECT 0.7000 246.6500 479.0000 246.9500 ;
      RECT 0.0000 244.9500 479.0000 246.6500 ;
      RECT 0.7000 244.6500 479.0000 244.9500 ;
      RECT 0.0000 242.9500 479.0000 244.6500 ;
      RECT 0.7000 242.6500 479.0000 242.9500 ;
      RECT 0.0000 240.9500 479.0000 242.6500 ;
      RECT 0.7000 240.6500 479.0000 240.9500 ;
      RECT 0.0000 238.9500 479.0000 240.6500 ;
      RECT 0.7000 238.6500 479.0000 238.9500 ;
      RECT 0.0000 236.9500 479.0000 238.6500 ;
      RECT 0.7000 236.6500 479.0000 236.9500 ;
      RECT 0.0000 234.9500 479.0000 236.6500 ;
      RECT 0.7000 234.6500 479.0000 234.9500 ;
      RECT 0.0000 232.9500 479.0000 234.6500 ;
      RECT 0.7000 232.6500 479.0000 232.9500 ;
      RECT 0.0000 230.9500 479.0000 232.6500 ;
      RECT 0.7000 230.6500 479.0000 230.9500 ;
      RECT 0.0000 228.9500 479.0000 230.6500 ;
      RECT 0.7000 228.6500 479.0000 228.9500 ;
      RECT 0.0000 226.9500 479.0000 228.6500 ;
      RECT 0.7000 226.6500 479.0000 226.9500 ;
      RECT 0.0000 224.9500 479.0000 226.6500 ;
      RECT 0.7000 224.6500 479.0000 224.9500 ;
      RECT 0.0000 222.9500 479.0000 224.6500 ;
      RECT 0.7000 222.6500 479.0000 222.9500 ;
      RECT 0.0000 220.9500 479.0000 222.6500 ;
      RECT 0.7000 220.6500 479.0000 220.9500 ;
      RECT 0.0000 218.9500 479.0000 220.6500 ;
      RECT 0.7000 218.6500 479.0000 218.9500 ;
      RECT 0.0000 216.9500 479.0000 218.6500 ;
      RECT 0.7000 216.6500 479.0000 216.9500 ;
      RECT 0.0000 214.9500 479.0000 216.6500 ;
      RECT 0.7000 214.6500 479.0000 214.9500 ;
      RECT 0.0000 212.9500 479.0000 214.6500 ;
      RECT 0.7000 212.6500 479.0000 212.9500 ;
      RECT 0.0000 210.9500 479.0000 212.6500 ;
      RECT 0.7000 210.6500 479.0000 210.9500 ;
      RECT 0.0000 208.9500 479.0000 210.6500 ;
      RECT 0.7000 208.6500 479.0000 208.9500 ;
      RECT 0.0000 206.9500 479.0000 208.6500 ;
      RECT 0.7000 206.6500 479.0000 206.9500 ;
      RECT 0.0000 204.9500 479.0000 206.6500 ;
      RECT 0.7000 204.6500 479.0000 204.9500 ;
      RECT 0.0000 202.9500 479.0000 204.6500 ;
      RECT 0.7000 202.6500 479.0000 202.9500 ;
      RECT 0.0000 200.9500 479.0000 202.6500 ;
      RECT 0.7000 200.6500 479.0000 200.9500 ;
      RECT 0.0000 198.9500 479.0000 200.6500 ;
      RECT 0.7000 198.6500 479.0000 198.9500 ;
      RECT 0.0000 196.9500 479.0000 198.6500 ;
      RECT 0.7000 196.6500 479.0000 196.9500 ;
      RECT 0.0000 194.9500 479.0000 196.6500 ;
      RECT 0.7000 194.6500 479.0000 194.9500 ;
      RECT 0.0000 192.9500 479.0000 194.6500 ;
      RECT 0.7000 192.6500 479.0000 192.9500 ;
      RECT 0.0000 190.9500 479.0000 192.6500 ;
      RECT 0.7000 190.6500 479.0000 190.9500 ;
      RECT 0.0000 188.9500 479.0000 190.6500 ;
      RECT 0.7000 188.6500 479.0000 188.9500 ;
      RECT 0.0000 186.9500 479.0000 188.6500 ;
      RECT 0.7000 186.6500 479.0000 186.9500 ;
      RECT 0.0000 184.9500 479.0000 186.6500 ;
      RECT 0.7000 184.6500 479.0000 184.9500 ;
      RECT 0.0000 182.9500 479.0000 184.6500 ;
      RECT 0.7000 182.6500 479.0000 182.9500 ;
      RECT 0.0000 180.9500 479.0000 182.6500 ;
      RECT 0.7000 180.6500 479.0000 180.9500 ;
      RECT 0.0000 178.9500 479.0000 180.6500 ;
      RECT 0.7000 178.6500 479.0000 178.9500 ;
      RECT 0.0000 176.9500 479.0000 178.6500 ;
      RECT 0.7000 176.6500 479.0000 176.9500 ;
      RECT 0.0000 174.9500 479.0000 176.6500 ;
      RECT 0.7000 174.6500 479.0000 174.9500 ;
      RECT 0.0000 172.9500 479.0000 174.6500 ;
      RECT 0.7000 172.6500 479.0000 172.9500 ;
      RECT 0.0000 170.9500 479.0000 172.6500 ;
      RECT 0.7000 170.6500 479.0000 170.9500 ;
      RECT 0.0000 168.9500 479.0000 170.6500 ;
      RECT 0.7000 168.6500 479.0000 168.9500 ;
      RECT 0.0000 166.9500 479.0000 168.6500 ;
      RECT 0.7000 166.6500 479.0000 166.9500 ;
      RECT 0.0000 164.9500 479.0000 166.6500 ;
      RECT 0.7000 164.6500 479.0000 164.9500 ;
      RECT 0.0000 162.9500 479.0000 164.6500 ;
      RECT 0.7000 162.6500 479.0000 162.9500 ;
      RECT 0.0000 160.9500 479.0000 162.6500 ;
      RECT 0.7000 160.6500 479.0000 160.9500 ;
      RECT 0.0000 158.9500 479.0000 160.6500 ;
      RECT 0.7000 158.6500 479.0000 158.9500 ;
      RECT 0.0000 156.9500 479.0000 158.6500 ;
      RECT 0.7000 156.6500 479.0000 156.9500 ;
      RECT 0.0000 0.7600 479.0000 156.6500 ;
      RECT 399.5100 0.0000 479.0000 0.7600 ;
      RECT 398.5100 0.0000 399.0900 0.7600 ;
      RECT 397.5100 0.0000 398.0900 0.7600 ;
      RECT 396.5100 0.0000 397.0900 0.7600 ;
      RECT 395.5100 0.0000 396.0900 0.7600 ;
      RECT 394.5100 0.0000 395.0900 0.7600 ;
      RECT 393.5100 0.0000 394.0900 0.7600 ;
      RECT 392.5100 0.0000 393.0900 0.7600 ;
      RECT 391.5100 0.0000 392.0900 0.7600 ;
      RECT 390.5100 0.0000 391.0900 0.7600 ;
      RECT 389.5100 0.0000 390.0900 0.7600 ;
      RECT 388.5100 0.0000 389.0900 0.7600 ;
      RECT 387.5100 0.0000 388.0900 0.7600 ;
      RECT 386.5100 0.0000 387.0900 0.7600 ;
      RECT 385.5100 0.0000 386.0900 0.7600 ;
      RECT 384.5100 0.0000 385.0900 0.7600 ;
      RECT 383.5100 0.0000 384.0900 0.7600 ;
      RECT 382.5100 0.0000 383.0900 0.7600 ;
      RECT 381.5100 0.0000 382.0900 0.7600 ;
      RECT 380.5100 0.0000 381.0900 0.7600 ;
      RECT 379.5100 0.0000 380.0900 0.7600 ;
      RECT 378.5100 0.0000 379.0900 0.7600 ;
      RECT 377.5100 0.0000 378.0900 0.7600 ;
      RECT 376.5100 0.0000 377.0900 0.7600 ;
      RECT 375.5100 0.0000 376.0900 0.7600 ;
      RECT 374.5100 0.0000 375.0900 0.7600 ;
      RECT 373.5100 0.0000 374.0900 0.7600 ;
      RECT 372.5100 0.0000 373.0900 0.7600 ;
      RECT 371.5100 0.0000 372.0900 0.7600 ;
      RECT 370.5100 0.0000 371.0900 0.7600 ;
      RECT 369.5100 0.0000 370.0900 0.7600 ;
      RECT 368.5100 0.0000 369.0900 0.7600 ;
      RECT 367.5100 0.0000 368.0900 0.7600 ;
      RECT 366.5100 0.0000 367.0900 0.7600 ;
      RECT 365.5100 0.0000 366.0900 0.7600 ;
      RECT 364.5100 0.0000 365.0900 0.7600 ;
      RECT 363.5100 0.0000 364.0900 0.7600 ;
      RECT 362.5100 0.0000 363.0900 0.7600 ;
      RECT 361.5100 0.0000 362.0900 0.7600 ;
      RECT 360.5100 0.0000 361.0900 0.7600 ;
      RECT 359.5100 0.0000 360.0900 0.7600 ;
      RECT 358.5100 0.0000 359.0900 0.7600 ;
      RECT 357.5100 0.0000 358.0900 0.7600 ;
      RECT 356.5100 0.0000 357.0900 0.7600 ;
      RECT 355.5100 0.0000 356.0900 0.7600 ;
      RECT 354.5100 0.0000 355.0900 0.7600 ;
      RECT 353.5100 0.0000 354.0900 0.7600 ;
      RECT 352.5100 0.0000 353.0900 0.7600 ;
      RECT 351.5100 0.0000 352.0900 0.7600 ;
      RECT 350.5100 0.0000 351.0900 0.7600 ;
      RECT 349.5100 0.0000 350.0900 0.7600 ;
      RECT 348.5100 0.0000 349.0900 0.7600 ;
      RECT 347.5100 0.0000 348.0900 0.7600 ;
      RECT 346.5100 0.0000 347.0900 0.7600 ;
      RECT 345.5100 0.0000 346.0900 0.7600 ;
      RECT 344.5100 0.0000 345.0900 0.7600 ;
      RECT 343.5100 0.0000 344.0900 0.7600 ;
      RECT 342.5100 0.0000 343.0900 0.7600 ;
      RECT 341.5100 0.0000 342.0900 0.7600 ;
      RECT 340.5100 0.0000 341.0900 0.7600 ;
      RECT 339.5100 0.0000 340.0900 0.7600 ;
      RECT 338.5100 0.0000 339.0900 0.7600 ;
      RECT 337.5100 0.0000 338.0900 0.7600 ;
      RECT 336.5100 0.0000 337.0900 0.7600 ;
      RECT 335.5100 0.0000 336.0900 0.7600 ;
      RECT 334.5100 0.0000 335.0900 0.7600 ;
      RECT 333.5100 0.0000 334.0900 0.7600 ;
      RECT 332.5100 0.0000 333.0900 0.7600 ;
      RECT 331.5100 0.0000 332.0900 0.7600 ;
      RECT 330.5100 0.0000 331.0900 0.7600 ;
      RECT 329.5100 0.0000 330.0900 0.7600 ;
      RECT 328.5100 0.0000 329.0900 0.7600 ;
      RECT 327.5100 0.0000 328.0900 0.7600 ;
      RECT 326.5100 0.0000 327.0900 0.7600 ;
      RECT 325.5100 0.0000 326.0900 0.7600 ;
      RECT 324.5100 0.0000 325.0900 0.7600 ;
      RECT 323.5100 0.0000 324.0900 0.7600 ;
      RECT 322.5100 0.0000 323.0900 0.7600 ;
      RECT 321.5100 0.0000 322.0900 0.7600 ;
      RECT 320.5100 0.0000 321.0900 0.7600 ;
      RECT 319.5100 0.0000 320.0900 0.7600 ;
      RECT 318.5100 0.0000 319.0900 0.7600 ;
      RECT 317.5100 0.0000 318.0900 0.7600 ;
      RECT 316.5100 0.0000 317.0900 0.7600 ;
      RECT 315.5100 0.0000 316.0900 0.7600 ;
      RECT 314.5100 0.0000 315.0900 0.7600 ;
      RECT 313.5100 0.0000 314.0900 0.7600 ;
      RECT 312.5100 0.0000 313.0900 0.7600 ;
      RECT 311.5100 0.0000 312.0900 0.7600 ;
      RECT 310.5100 0.0000 311.0900 0.7600 ;
      RECT 309.5100 0.0000 310.0900 0.7600 ;
      RECT 308.5100 0.0000 309.0900 0.7600 ;
      RECT 307.5100 0.0000 308.0900 0.7600 ;
      RECT 306.5100 0.0000 307.0900 0.7600 ;
      RECT 305.5100 0.0000 306.0900 0.7600 ;
      RECT 304.5100 0.0000 305.0900 0.7600 ;
      RECT 303.5100 0.0000 304.0900 0.7600 ;
      RECT 302.5100 0.0000 303.0900 0.7600 ;
      RECT 301.5100 0.0000 302.0900 0.7600 ;
      RECT 300.5100 0.0000 301.0900 0.7600 ;
      RECT 299.5100 0.0000 300.0900 0.7600 ;
      RECT 298.5100 0.0000 299.0900 0.7600 ;
      RECT 297.5100 0.0000 298.0900 0.7600 ;
      RECT 296.5100 0.0000 297.0900 0.7600 ;
      RECT 295.5100 0.0000 296.0900 0.7600 ;
      RECT 294.5100 0.0000 295.0900 0.7600 ;
      RECT 293.5100 0.0000 294.0900 0.7600 ;
      RECT 292.5100 0.0000 293.0900 0.7600 ;
      RECT 291.5100 0.0000 292.0900 0.7600 ;
      RECT 290.5100 0.0000 291.0900 0.7600 ;
      RECT 289.5100 0.0000 290.0900 0.7600 ;
      RECT 288.5100 0.0000 289.0900 0.7600 ;
      RECT 287.5100 0.0000 288.0900 0.7600 ;
      RECT 286.5100 0.0000 287.0900 0.7600 ;
      RECT 285.5100 0.0000 286.0900 0.7600 ;
      RECT 284.5100 0.0000 285.0900 0.7600 ;
      RECT 283.5100 0.0000 284.0900 0.7600 ;
      RECT 282.5100 0.0000 283.0900 0.7600 ;
      RECT 281.5100 0.0000 282.0900 0.7600 ;
      RECT 280.5100 0.0000 281.0900 0.7600 ;
      RECT 279.5100 0.0000 280.0900 0.7600 ;
      RECT 278.5100 0.0000 279.0900 0.7600 ;
      RECT 277.5100 0.0000 278.0900 0.7600 ;
      RECT 276.5100 0.0000 277.0900 0.7600 ;
      RECT 275.5100 0.0000 276.0900 0.7600 ;
      RECT 274.5100 0.0000 275.0900 0.7600 ;
      RECT 273.5100 0.0000 274.0900 0.7600 ;
      RECT 272.5100 0.0000 273.0900 0.7600 ;
      RECT 271.5100 0.0000 272.0900 0.7600 ;
      RECT 270.5100 0.0000 271.0900 0.7600 ;
      RECT 269.5100 0.0000 270.0900 0.7600 ;
      RECT 268.5100 0.0000 269.0900 0.7600 ;
      RECT 267.5100 0.0000 268.0900 0.7600 ;
      RECT 266.5100 0.0000 267.0900 0.7600 ;
      RECT 265.5100 0.0000 266.0900 0.7600 ;
      RECT 264.5100 0.0000 265.0900 0.7600 ;
      RECT 263.5100 0.0000 264.0900 0.7600 ;
      RECT 262.5100 0.0000 263.0900 0.7600 ;
      RECT 261.5100 0.0000 262.0900 0.7600 ;
      RECT 260.5100 0.0000 261.0900 0.7600 ;
      RECT 259.5100 0.0000 260.0900 0.7600 ;
      RECT 258.5100 0.0000 259.0900 0.7600 ;
      RECT 257.5100 0.0000 258.0900 0.7600 ;
      RECT 256.5100 0.0000 257.0900 0.7600 ;
      RECT 255.5100 0.0000 256.0900 0.7600 ;
      RECT 254.5100 0.0000 255.0900 0.7600 ;
      RECT 253.5100 0.0000 254.0900 0.7600 ;
      RECT 252.5100 0.0000 253.0900 0.7600 ;
      RECT 251.5100 0.0000 252.0900 0.7600 ;
      RECT 250.5100 0.0000 251.0900 0.7600 ;
      RECT 249.5100 0.0000 250.0900 0.7600 ;
      RECT 248.5100 0.0000 249.0900 0.7600 ;
      RECT 247.5100 0.0000 248.0900 0.7600 ;
      RECT 246.5100 0.0000 247.0900 0.7600 ;
      RECT 245.5100 0.0000 246.0900 0.7600 ;
      RECT 244.5100 0.0000 245.0900 0.7600 ;
      RECT 243.5100 0.0000 244.0900 0.7600 ;
      RECT 242.5100 0.0000 243.0900 0.7600 ;
      RECT 241.5100 0.0000 242.0900 0.7600 ;
      RECT 240.5100 0.0000 241.0900 0.7600 ;
      RECT 239.5100 0.0000 240.0900 0.7600 ;
      RECT 238.5100 0.0000 239.0900 0.7600 ;
      RECT 237.5100 0.0000 238.0900 0.7600 ;
      RECT 236.5100 0.0000 237.0900 0.7600 ;
      RECT 235.5100 0.0000 236.0900 0.7600 ;
      RECT 234.5100 0.0000 235.0900 0.7600 ;
      RECT 233.5100 0.0000 234.0900 0.7600 ;
      RECT 232.5100 0.0000 233.0900 0.7600 ;
      RECT 231.5100 0.0000 232.0900 0.7600 ;
      RECT 230.5100 0.0000 231.0900 0.7600 ;
      RECT 229.5100 0.0000 230.0900 0.7600 ;
      RECT 228.5100 0.0000 229.0900 0.7600 ;
      RECT 227.5100 0.0000 228.0900 0.7600 ;
      RECT 226.5100 0.0000 227.0900 0.7600 ;
      RECT 225.5100 0.0000 226.0900 0.7600 ;
      RECT 224.5100 0.0000 225.0900 0.7600 ;
      RECT 223.5100 0.0000 224.0900 0.7600 ;
      RECT 222.5100 0.0000 223.0900 0.7600 ;
      RECT 221.5100 0.0000 222.0900 0.7600 ;
      RECT 220.5100 0.0000 221.0900 0.7600 ;
      RECT 219.5100 0.0000 220.0900 0.7600 ;
      RECT 218.5100 0.0000 219.0900 0.7600 ;
      RECT 217.5100 0.0000 218.0900 0.7600 ;
      RECT 216.5100 0.0000 217.0900 0.7600 ;
      RECT 215.5100 0.0000 216.0900 0.7600 ;
      RECT 214.5100 0.0000 215.0900 0.7600 ;
      RECT 213.5100 0.0000 214.0900 0.7600 ;
      RECT 212.5100 0.0000 213.0900 0.7600 ;
      RECT 211.5100 0.0000 212.0900 0.7600 ;
      RECT 210.5100 0.0000 211.0900 0.7600 ;
      RECT 209.5100 0.0000 210.0900 0.7600 ;
      RECT 208.5100 0.0000 209.0900 0.7600 ;
      RECT 207.5100 0.0000 208.0900 0.7600 ;
      RECT 206.5100 0.0000 207.0900 0.7600 ;
      RECT 205.5100 0.0000 206.0900 0.7600 ;
      RECT 204.5100 0.0000 205.0900 0.7600 ;
      RECT 203.5100 0.0000 204.0900 0.7600 ;
      RECT 202.5100 0.0000 203.0900 0.7600 ;
      RECT 201.5100 0.0000 202.0900 0.7600 ;
      RECT 200.5100 0.0000 201.0900 0.7600 ;
      RECT 199.5100 0.0000 200.0900 0.7600 ;
      RECT 198.5100 0.0000 199.0900 0.7600 ;
      RECT 197.5100 0.0000 198.0900 0.7600 ;
      RECT 196.5100 0.0000 197.0900 0.7600 ;
      RECT 195.5100 0.0000 196.0900 0.7600 ;
      RECT 194.5100 0.0000 195.0900 0.7600 ;
      RECT 193.5100 0.0000 194.0900 0.7600 ;
      RECT 192.5100 0.0000 193.0900 0.7600 ;
      RECT 191.5100 0.0000 192.0900 0.7600 ;
      RECT 190.5100 0.0000 191.0900 0.7600 ;
      RECT 189.5100 0.0000 190.0900 0.7600 ;
      RECT 188.5100 0.0000 189.0900 0.7600 ;
      RECT 187.5100 0.0000 188.0900 0.7600 ;
      RECT 186.5100 0.0000 187.0900 0.7600 ;
      RECT 185.5100 0.0000 186.0900 0.7600 ;
      RECT 184.5100 0.0000 185.0900 0.7600 ;
      RECT 183.5100 0.0000 184.0900 0.7600 ;
      RECT 182.5100 0.0000 183.0900 0.7600 ;
      RECT 181.5100 0.0000 182.0900 0.7600 ;
      RECT 180.5100 0.0000 181.0900 0.7600 ;
      RECT 179.5100 0.0000 180.0900 0.7600 ;
      RECT 178.5100 0.0000 179.0900 0.7600 ;
      RECT 177.5100 0.0000 178.0900 0.7600 ;
      RECT 176.5100 0.0000 177.0900 0.7600 ;
      RECT 175.5100 0.0000 176.0900 0.7600 ;
      RECT 174.5100 0.0000 175.0900 0.7600 ;
      RECT 173.5100 0.0000 174.0900 0.7600 ;
      RECT 172.5100 0.0000 173.0900 0.7600 ;
      RECT 171.5100 0.0000 172.0900 0.7600 ;
      RECT 170.5100 0.0000 171.0900 0.7600 ;
      RECT 169.5100 0.0000 170.0900 0.7600 ;
      RECT 168.5100 0.0000 169.0900 0.7600 ;
      RECT 167.5100 0.0000 168.0900 0.7600 ;
      RECT 166.5100 0.0000 167.0900 0.7600 ;
      RECT 165.5100 0.0000 166.0900 0.7600 ;
      RECT 164.5100 0.0000 165.0900 0.7600 ;
      RECT 163.5100 0.0000 164.0900 0.7600 ;
      RECT 162.5100 0.0000 163.0900 0.7600 ;
      RECT 161.5100 0.0000 162.0900 0.7600 ;
      RECT 160.5100 0.0000 161.0900 0.7600 ;
      RECT 159.5100 0.0000 160.0900 0.7600 ;
      RECT 158.5100 0.0000 159.0900 0.7600 ;
      RECT 157.5100 0.0000 158.0900 0.7600 ;
      RECT 156.5100 0.0000 157.0900 0.7600 ;
      RECT 155.5100 0.0000 156.0900 0.7600 ;
      RECT 154.5100 0.0000 155.0900 0.7600 ;
      RECT 153.5100 0.0000 154.0900 0.7600 ;
      RECT 152.5100 0.0000 153.0900 0.7600 ;
      RECT 151.5100 0.0000 152.0900 0.7600 ;
      RECT 150.5100 0.0000 151.0900 0.7600 ;
      RECT 149.5100 0.0000 150.0900 0.7600 ;
      RECT 148.5100 0.0000 149.0900 0.7600 ;
      RECT 147.5100 0.0000 148.0900 0.7600 ;
      RECT 146.5100 0.0000 147.0900 0.7600 ;
      RECT 145.5100 0.0000 146.0900 0.7600 ;
      RECT 144.5100 0.0000 145.0900 0.7600 ;
      RECT 143.5100 0.0000 144.0900 0.7600 ;
      RECT 142.5100 0.0000 143.0900 0.7600 ;
      RECT 141.5100 0.0000 142.0900 0.7600 ;
      RECT 140.5100 0.0000 141.0900 0.7600 ;
      RECT 139.5100 0.0000 140.0900 0.7600 ;
      RECT 138.5100 0.0000 139.0900 0.7600 ;
      RECT 137.5100 0.0000 138.0900 0.7600 ;
      RECT 136.5100 0.0000 137.0900 0.7600 ;
      RECT 135.5100 0.0000 136.0900 0.7600 ;
      RECT 134.5100 0.0000 135.0900 0.7600 ;
      RECT 133.5100 0.0000 134.0900 0.7600 ;
      RECT 132.5100 0.0000 133.0900 0.7600 ;
      RECT 131.5100 0.0000 132.0900 0.7600 ;
      RECT 130.5100 0.0000 131.0900 0.7600 ;
      RECT 129.5100 0.0000 130.0900 0.7600 ;
      RECT 128.5100 0.0000 129.0900 0.7600 ;
      RECT 127.5100 0.0000 128.0900 0.7600 ;
      RECT 126.5100 0.0000 127.0900 0.7600 ;
      RECT 125.5100 0.0000 126.0900 0.7600 ;
      RECT 124.5100 0.0000 125.0900 0.7600 ;
      RECT 123.5100 0.0000 124.0900 0.7600 ;
      RECT 122.5100 0.0000 123.0900 0.7600 ;
      RECT 121.5100 0.0000 122.0900 0.7600 ;
      RECT 120.5100 0.0000 121.0900 0.7600 ;
      RECT 119.5100 0.0000 120.0900 0.7600 ;
      RECT 118.5100 0.0000 119.0900 0.7600 ;
      RECT 117.5100 0.0000 118.0900 0.7600 ;
      RECT 116.5100 0.0000 117.0900 0.7600 ;
      RECT 115.5100 0.0000 116.0900 0.7600 ;
      RECT 114.5100 0.0000 115.0900 0.7600 ;
      RECT 113.5100 0.0000 114.0900 0.7600 ;
      RECT 112.5100 0.0000 113.0900 0.7600 ;
      RECT 111.5100 0.0000 112.0900 0.7600 ;
      RECT 110.5100 0.0000 111.0900 0.7600 ;
      RECT 109.5100 0.0000 110.0900 0.7600 ;
      RECT 108.5100 0.0000 109.0900 0.7600 ;
      RECT 107.5100 0.0000 108.0900 0.7600 ;
      RECT 106.5100 0.0000 107.0900 0.7600 ;
      RECT 105.5100 0.0000 106.0900 0.7600 ;
      RECT 104.5100 0.0000 105.0900 0.7600 ;
      RECT 103.5100 0.0000 104.0900 0.7600 ;
      RECT 102.5100 0.0000 103.0900 0.7600 ;
      RECT 101.5100 0.0000 102.0900 0.7600 ;
      RECT 100.5100 0.0000 101.0900 0.7600 ;
      RECT 99.5100 0.0000 100.0900 0.7600 ;
      RECT 98.5100 0.0000 99.0900 0.7600 ;
      RECT 97.5100 0.0000 98.0900 0.7600 ;
      RECT 96.5100 0.0000 97.0900 0.7600 ;
      RECT 95.5100 0.0000 96.0900 0.7600 ;
      RECT 94.5100 0.0000 95.0900 0.7600 ;
      RECT 93.5100 0.0000 94.0900 0.7600 ;
      RECT 92.5100 0.0000 93.0900 0.7600 ;
      RECT 91.5100 0.0000 92.0900 0.7600 ;
      RECT 90.5100 0.0000 91.0900 0.7600 ;
      RECT 89.5100 0.0000 90.0900 0.7600 ;
      RECT 88.5100 0.0000 89.0900 0.7600 ;
      RECT 87.5100 0.0000 88.0900 0.7600 ;
      RECT 86.5100 0.0000 87.0900 0.7600 ;
      RECT 85.5100 0.0000 86.0900 0.7600 ;
      RECT 84.5100 0.0000 85.0900 0.7600 ;
      RECT 83.5100 0.0000 84.0900 0.7600 ;
      RECT 82.5100 0.0000 83.0900 0.7600 ;
      RECT 81.5100 0.0000 82.0900 0.7600 ;
      RECT 80.5100 0.0000 81.0900 0.7600 ;
      RECT 0.0000 0.0000 80.0900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 479.0000 477.2000 ;
  END
END core

END LIBRARY
