/home/linux/ieng6/ee260bwi25/b8kang/step3/sram/pnr/sram_w16.lef