##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sun Mar  9 15:37:23 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 438.8000 BY 437.6000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 200.5500 0.6000 200.6500 ;
    END
  END clk
  PIN sum_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 219.0500 0.0000 219.1500 0.6000 ;
    END
  END sum_out[159]
  PIN sum_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.2500 0.0000 218.3500 0.6000 ;
    END
  END sum_out[158]
  PIN sum_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.4500 0.0000 217.5500 0.6000 ;
    END
  END sum_out[157]
  PIN sum_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 216.6500 0.0000 216.7500 0.6000 ;
    END
  END sum_out[156]
  PIN sum_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.8500 0.0000 215.9500 0.6000 ;
    END
  END sum_out[155]
  PIN sum_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.0500 0.0000 215.1500 0.6000 ;
    END
  END sum_out[154]
  PIN sum_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 214.2500 0.0000 214.3500 0.6000 ;
    END
  END sum_out[153]
  PIN sum_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.4500 0.0000 213.5500 0.6000 ;
    END
  END sum_out[152]
  PIN sum_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.6500 0.0000 212.7500 0.6000 ;
    END
  END sum_out[151]
  PIN sum_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 211.8500 0.0000 211.9500 0.6000 ;
    END
  END sum_out[150]
  PIN sum_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 211.0500 0.0000 211.1500 0.6000 ;
    END
  END sum_out[149]
  PIN sum_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.2500 0.0000 210.3500 0.6000 ;
    END
  END sum_out[148]
  PIN sum_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.4500 0.0000 209.5500 0.6000 ;
    END
  END sum_out[147]
  PIN sum_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 208.6500 0.0000 208.7500 0.6000 ;
    END
  END sum_out[146]
  PIN sum_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.8500 0.0000 207.9500 0.6000 ;
    END
  END sum_out[145]
  PIN sum_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.0500 0.0000 207.1500 0.6000 ;
    END
  END sum_out[144]
  PIN sum_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 206.2500 0.0000 206.3500 0.6000 ;
    END
  END sum_out[143]
  PIN sum_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.4500 0.0000 205.5500 0.6000 ;
    END
  END sum_out[142]
  PIN sum_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.6500 0.0000 204.7500 0.6000 ;
    END
  END sum_out[141]
  PIN sum_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 203.8500 0.0000 203.9500 0.6000 ;
    END
  END sum_out[140]
  PIN sum_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 203.0500 0.0000 203.1500 0.6000 ;
    END
  END sum_out[139]
  PIN sum_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.2500 0.0000 202.3500 0.6000 ;
    END
  END sum_out[138]
  PIN sum_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.4500 0.0000 201.5500 0.6000 ;
    END
  END sum_out[137]
  PIN sum_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 200.6500 0.0000 200.7500 0.6000 ;
    END
  END sum_out[136]
  PIN sum_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.8500 0.0000 199.9500 0.6000 ;
    END
  END sum_out[135]
  PIN sum_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.0500 0.0000 199.1500 0.6000 ;
    END
  END sum_out[134]
  PIN sum_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 198.2500 0.0000 198.3500 0.6000 ;
    END
  END sum_out[133]
  PIN sum_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.4500 0.0000 197.5500 0.6000 ;
    END
  END sum_out[132]
  PIN sum_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.6500 0.0000 196.7500 0.6000 ;
    END
  END sum_out[131]
  PIN sum_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 195.8500 0.0000 195.9500 0.6000 ;
    END
  END sum_out[130]
  PIN sum_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 195.0500 0.0000 195.1500 0.6000 ;
    END
  END sum_out[129]
  PIN sum_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.2500 0.0000 194.3500 0.6000 ;
    END
  END sum_out[128]
  PIN sum_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.4500 0.0000 193.5500 0.6000 ;
    END
  END sum_out[127]
  PIN sum_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 192.6500 0.0000 192.7500 0.6000 ;
    END
  END sum_out[126]
  PIN sum_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.8500 0.0000 191.9500 0.6000 ;
    END
  END sum_out[125]
  PIN sum_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.0500 0.0000 191.1500 0.6000 ;
    END
  END sum_out[124]
  PIN sum_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 190.2500 0.0000 190.3500 0.6000 ;
    END
  END sum_out[123]
  PIN sum_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.4500 0.0000 189.5500 0.6000 ;
    END
  END sum_out[122]
  PIN sum_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.6500 0.0000 188.7500 0.6000 ;
    END
  END sum_out[121]
  PIN sum_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 187.8500 0.0000 187.9500 0.6000 ;
    END
  END sum_out[120]
  PIN sum_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 187.0500 0.0000 187.1500 0.6000 ;
    END
  END sum_out[119]
  PIN sum_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.2500 0.0000 186.3500 0.6000 ;
    END
  END sum_out[118]
  PIN sum_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.4500 0.0000 185.5500 0.6000 ;
    END
  END sum_out[117]
  PIN sum_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.6500 0.0000 184.7500 0.6000 ;
    END
  END sum_out[116]
  PIN sum_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.8500 0.0000 183.9500 0.6000 ;
    END
  END sum_out[115]
  PIN sum_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.0500 0.0000 183.1500 0.6000 ;
    END
  END sum_out[114]
  PIN sum_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.2500 0.0000 182.3500 0.6000 ;
    END
  END sum_out[113]
  PIN sum_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.4500 0.0000 181.5500 0.6000 ;
    END
  END sum_out[112]
  PIN sum_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.6500 0.0000 180.7500 0.6000 ;
    END
  END sum_out[111]
  PIN sum_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.8500 0.0000 179.9500 0.6000 ;
    END
  END sum_out[110]
  PIN sum_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.0500 0.0000 179.1500 0.6000 ;
    END
  END sum_out[109]
  PIN sum_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.2500 0.0000 178.3500 0.6000 ;
    END
  END sum_out[108]
  PIN sum_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.4500 0.0000 177.5500 0.6000 ;
    END
  END sum_out[107]
  PIN sum_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.6500 0.0000 176.7500 0.6000 ;
    END
  END sum_out[106]
  PIN sum_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.8500 0.0000 175.9500 0.6000 ;
    END
  END sum_out[105]
  PIN sum_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.0500 0.0000 175.1500 0.6000 ;
    END
  END sum_out[104]
  PIN sum_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.2500 0.0000 174.3500 0.6000 ;
    END
  END sum_out[103]
  PIN sum_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.4500 0.0000 173.5500 0.6000 ;
    END
  END sum_out[102]
  PIN sum_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.6500 0.0000 172.7500 0.6000 ;
    END
  END sum_out[101]
  PIN sum_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.8500 0.0000 171.9500 0.6000 ;
    END
  END sum_out[100]
  PIN sum_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.0500 0.0000 171.1500 0.6000 ;
    END
  END sum_out[99]
  PIN sum_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.2500 0.0000 170.3500 0.6000 ;
    END
  END sum_out[98]
  PIN sum_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.4500 0.0000 169.5500 0.6000 ;
    END
  END sum_out[97]
  PIN sum_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.6500 0.0000 168.7500 0.6000 ;
    END
  END sum_out[96]
  PIN sum_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.8500 0.0000 167.9500 0.6000 ;
    END
  END sum_out[95]
  PIN sum_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.0500 0.0000 167.1500 0.6000 ;
    END
  END sum_out[94]
  PIN sum_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.2500 0.0000 166.3500 0.6000 ;
    END
  END sum_out[93]
  PIN sum_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.4500 0.0000 165.5500 0.6000 ;
    END
  END sum_out[92]
  PIN sum_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.6500 0.0000 164.7500 0.6000 ;
    END
  END sum_out[91]
  PIN sum_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.8500 0.0000 163.9500 0.6000 ;
    END
  END sum_out[90]
  PIN sum_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.0500 0.0000 163.1500 0.6000 ;
    END
  END sum_out[89]
  PIN sum_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.2500 0.0000 162.3500 0.6000 ;
    END
  END sum_out[88]
  PIN sum_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.4500 0.0000 161.5500 0.6000 ;
    END
  END sum_out[87]
  PIN sum_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.6500 0.0000 160.7500 0.6000 ;
    END
  END sum_out[86]
  PIN sum_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.8500 0.0000 159.9500 0.6000 ;
    END
  END sum_out[85]
  PIN sum_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.0500 0.0000 159.1500 0.6000 ;
    END
  END sum_out[84]
  PIN sum_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.2500 0.0000 158.3500 0.6000 ;
    END
  END sum_out[83]
  PIN sum_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.4500 0.0000 157.5500 0.6000 ;
    END
  END sum_out[82]
  PIN sum_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.6500 0.0000 156.7500 0.6000 ;
    END
  END sum_out[81]
  PIN sum_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.8500 0.0000 155.9500 0.6000 ;
    END
  END sum_out[80]
  PIN sum_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.0500 0.0000 155.1500 0.6000 ;
    END
  END sum_out[79]
  PIN sum_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.2500 0.0000 154.3500 0.6000 ;
    END
  END sum_out[78]
  PIN sum_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.4500 0.0000 153.5500 0.6000 ;
    END
  END sum_out[77]
  PIN sum_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.6500 0.0000 152.7500 0.6000 ;
    END
  END sum_out[76]
  PIN sum_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.8500 0.0000 151.9500 0.6000 ;
    END
  END sum_out[75]
  PIN sum_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.0500 0.0000 151.1500 0.6000 ;
    END
  END sum_out[74]
  PIN sum_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.2500 0.0000 150.3500 0.6000 ;
    END
  END sum_out[73]
  PIN sum_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.4500 0.0000 149.5500 0.6000 ;
    END
  END sum_out[72]
  PIN sum_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.6500 0.0000 148.7500 0.6000 ;
    END
  END sum_out[71]
  PIN sum_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.8500 0.0000 147.9500 0.6000 ;
    END
  END sum_out[70]
  PIN sum_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.0500 0.0000 147.1500 0.6000 ;
    END
  END sum_out[69]
  PIN sum_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.2500 0.0000 146.3500 0.6000 ;
    END
  END sum_out[68]
  PIN sum_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.4500 0.0000 145.5500 0.6000 ;
    END
  END sum_out[67]
  PIN sum_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.6500 0.0000 144.7500 0.6000 ;
    END
  END sum_out[66]
  PIN sum_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.8500 0.0000 143.9500 0.6000 ;
    END
  END sum_out[65]
  PIN sum_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.0500 0.0000 143.1500 0.6000 ;
    END
  END sum_out[64]
  PIN sum_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 142.2500 0.0000 142.3500 0.6000 ;
    END
  END sum_out[63]
  PIN sum_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.4500 0.0000 141.5500 0.6000 ;
    END
  END sum_out[62]
  PIN sum_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.6500 0.0000 140.7500 0.6000 ;
    END
  END sum_out[61]
  PIN sum_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 139.8500 0.0000 139.9500 0.6000 ;
    END
  END sum_out[60]
  PIN sum_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 139.0500 0.0000 139.1500 0.6000 ;
    END
  END sum_out[59]
  PIN sum_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.2500 0.0000 138.3500 0.6000 ;
    END
  END sum_out[58]
  PIN sum_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.4500 0.0000 137.5500 0.6000 ;
    END
  END sum_out[57]
  PIN sum_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.6500 0.0000 136.7500 0.6000 ;
    END
  END sum_out[56]
  PIN sum_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.8500 0.0000 135.9500 0.6000 ;
    END
  END sum_out[55]
  PIN sum_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.0500 0.0000 135.1500 0.6000 ;
    END
  END sum_out[54]
  PIN sum_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.2500 0.0000 134.3500 0.6000 ;
    END
  END sum_out[53]
  PIN sum_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.4500 0.0000 133.5500 0.6000 ;
    END
  END sum_out[52]
  PIN sum_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.6500 0.0000 132.7500 0.6000 ;
    END
  END sum_out[51]
  PIN sum_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.8500 0.0000 131.9500 0.6000 ;
    END
  END sum_out[50]
  PIN sum_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.0500 0.0000 131.1500 0.6000 ;
    END
  END sum_out[49]
  PIN sum_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.2500 0.0000 130.3500 0.6000 ;
    END
  END sum_out[48]
  PIN sum_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.4500 0.0000 129.5500 0.6000 ;
    END
  END sum_out[47]
  PIN sum_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.6500 0.0000 128.7500 0.6000 ;
    END
  END sum_out[46]
  PIN sum_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.8500 0.0000 127.9500 0.6000 ;
    END
  END sum_out[45]
  PIN sum_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.0500 0.0000 127.1500 0.6000 ;
    END
  END sum_out[44]
  PIN sum_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 126.2500 0.0000 126.3500 0.6000 ;
    END
  END sum_out[43]
  PIN sum_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.4500 0.0000 125.5500 0.6000 ;
    END
  END sum_out[42]
  PIN sum_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.6500 0.0000 124.7500 0.6000 ;
    END
  END sum_out[41]
  PIN sum_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.8500 0.0000 123.9500 0.6000 ;
    END
  END sum_out[40]
  PIN sum_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.0500 0.0000 123.1500 0.6000 ;
    END
  END sum_out[39]
  PIN sum_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.2500 0.0000 122.3500 0.6000 ;
    END
  END sum_out[38]
  PIN sum_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.4500 0.0000 121.5500 0.6000 ;
    END
  END sum_out[37]
  PIN sum_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.6500 0.0000 120.7500 0.6000 ;
    END
  END sum_out[36]
  PIN sum_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.8500 0.0000 119.9500 0.6000 ;
    END
  END sum_out[35]
  PIN sum_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.0500 0.0000 119.1500 0.6000 ;
    END
  END sum_out[34]
  PIN sum_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 118.2500 0.0000 118.3500 0.6000 ;
    END
  END sum_out[33]
  PIN sum_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.4500 0.0000 117.5500 0.6000 ;
    END
  END sum_out[32]
  PIN sum_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.6500 0.0000 116.7500 0.6000 ;
    END
  END sum_out[31]
  PIN sum_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.8500 0.0000 115.9500 0.6000 ;
    END
  END sum_out[30]
  PIN sum_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.0500 0.0000 115.1500 0.6000 ;
    END
  END sum_out[29]
  PIN sum_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.2500 0.0000 114.3500 0.6000 ;
    END
  END sum_out[28]
  PIN sum_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.4500 0.0000 113.5500 0.6000 ;
    END
  END sum_out[27]
  PIN sum_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.6500 0.0000 112.7500 0.6000 ;
    END
  END sum_out[26]
  PIN sum_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.8500 0.0000 111.9500 0.6000 ;
    END
  END sum_out[25]
  PIN sum_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.0500 0.0000 111.1500 0.6000 ;
    END
  END sum_out[24]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 110.2500 0.0000 110.3500 0.6000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.4500 0.0000 109.5500 0.6000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.6500 0.0000 108.7500 0.6000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 107.8500 0.0000 107.9500 0.6000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 107.0500 0.0000 107.1500 0.6000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.2500 0.0000 106.3500 0.6000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.4500 0.0000 105.5500 0.6000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.6500 0.0000 104.7500 0.6000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.8500 0.0000 103.9500 0.6000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.0500 0.0000 103.1500 0.6000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 102.2500 0.0000 102.3500 0.6000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.4500 0.0000 101.5500 0.6000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.6500 0.0000 100.7500 0.6000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 99.8500 0.0000 99.9500 0.6000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 99.0500 0.0000 99.1500 0.6000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.2500 0.0000 98.3500 0.6000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.4500 0.0000 97.5500 0.6000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.6500 0.0000 96.7500 0.6000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.8500 0.0000 95.9500 0.6000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.0500 0.0000 95.1500 0.6000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 94.2500 0.0000 94.3500 0.6000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.4500 0.0000 93.5500 0.6000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.6500 0.0000 92.7500 0.6000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.8500 0.0000 91.9500 0.6000 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 251.7500 0.6000 251.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 250.9500 0.6000 251.0500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 250.1500 0.6000 250.2500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 249.3500 0.6000 249.4500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 248.5500 0.6000 248.6500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 247.7500 0.6000 247.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 246.9500 0.6000 247.0500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 246.1500 0.6000 246.2500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 245.3500 0.6000 245.4500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 244.5500 0.6000 244.6500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 243.7500 0.6000 243.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 242.9500 0.6000 243.0500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 242.1500 0.6000 242.2500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 241.3500 0.6000 241.4500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 240.5500 0.6000 240.6500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 239.7500 0.6000 239.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 238.9500 0.6000 239.0500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 238.1500 0.6000 238.2500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 237.3500 0.6000 237.4500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 236.5500 0.6000 236.6500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 235.7500 0.6000 235.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 234.9500 0.6000 235.0500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 234.1500 0.6000 234.2500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 233.3500 0.6000 233.4500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 232.5500 0.6000 232.6500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 231.7500 0.6000 231.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 230.9500 0.6000 231.0500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 230.1500 0.6000 230.2500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 229.3500 0.6000 229.4500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 228.5500 0.6000 228.6500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 227.7500 0.6000 227.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 226.9500 0.6000 227.0500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 226.1500 0.6000 226.2500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 225.3500 0.6000 225.4500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 224.5500 0.6000 224.6500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 223.7500 0.6000 223.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 222.9500 0.6000 223.0500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 222.1500 0.6000 222.2500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 221.3500 0.6000 221.4500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 220.5500 0.6000 220.6500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 219.7500 0.6000 219.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 218.9500 0.6000 219.0500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 218.1500 0.6000 218.2500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 217.3500 0.6000 217.4500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 216.5500 0.6000 216.6500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.7500 0.6000 215.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 214.9500 0.6000 215.0500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 214.1500 0.6000 214.2500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.3500 0.6000 213.4500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 212.5500 0.6000 212.6500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 211.7500 0.6000 211.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.9500 0.6000 211.0500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.1500 0.6000 210.2500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.3500 0.6000 209.4500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 208.5500 0.6000 208.6500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 207.7500 0.6000 207.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 206.9500 0.6000 207.0500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 206.1500 0.6000 206.2500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.3500 0.6000 205.4500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 204.5500 0.6000 204.6500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 203.7500 0.6000 203.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 202.9500 0.6000 203.0500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 202.1500 0.6000 202.2500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 201.3500 0.6000 201.4500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 347.0500 0.0000 347.1500 0.6000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.2500 0.0000 346.3500 0.6000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.4500 0.0000 345.5500 0.6000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 344.6500 0.0000 344.7500 0.6000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.8500 0.0000 343.9500 0.6000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.0500 0.0000 343.1500 0.6000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.2500 0.0000 342.3500 0.6000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.4500 0.0000 341.5500 0.6000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.6500 0.0000 340.7500 0.6000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.8500 0.0000 339.9500 0.6000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.0500 0.0000 339.1500 0.6000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.2500 0.0000 338.3500 0.6000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.4500 0.0000 337.5500 0.6000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.6500 0.0000 336.7500 0.6000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.8500 0.0000 335.9500 0.6000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.0500 0.0000 335.1500 0.6000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.2500 0.0000 334.3500 0.6000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.4500 0.0000 333.5500 0.6000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.6500 0.0000 332.7500 0.6000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.8500 0.0000 331.9500 0.6000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.0500 0.0000 331.1500 0.6000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.2500 0.0000 330.3500 0.6000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.4500 0.0000 329.5500 0.6000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 328.6500 0.0000 328.7500 0.6000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.8500 0.0000 327.9500 0.6000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.0500 0.0000 327.1500 0.6000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 326.2500 0.0000 326.3500 0.6000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.4500 0.0000 325.5500 0.6000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.6500 0.0000 324.7500 0.6000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.8500 0.0000 323.9500 0.6000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.0500 0.0000 323.1500 0.6000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.2500 0.0000 322.3500 0.6000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.4500 0.0000 321.5500 0.6000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 320.6500 0.0000 320.7500 0.6000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.8500 0.0000 319.9500 0.6000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.0500 0.0000 319.1500 0.6000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.2500 0.0000 318.3500 0.6000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.4500 0.0000 317.5500 0.6000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.6500 0.0000 316.7500 0.6000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.8500 0.0000 315.9500 0.6000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.0500 0.0000 315.1500 0.6000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.2500 0.0000 314.3500 0.6000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.4500 0.0000 313.5500 0.6000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.6500 0.0000 312.7500 0.6000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.8500 0.0000 311.9500 0.6000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.0500 0.0000 311.1500 0.6000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.2500 0.0000 310.3500 0.6000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.4500 0.0000 309.5500 0.6000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.6500 0.0000 308.7500 0.6000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.8500 0.0000 307.9500 0.6000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.0500 0.0000 307.1500 0.6000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.2500 0.0000 306.3500 0.6000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.4500 0.0000 305.5500 0.6000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 304.6500 0.0000 304.7500 0.6000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.8500 0.0000 303.9500 0.6000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.0500 0.0000 303.1500 0.6000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 302.2500 0.0000 302.3500 0.6000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.4500 0.0000 301.5500 0.6000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.6500 0.0000 300.7500 0.6000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.8500 0.0000 299.9500 0.6000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.0500 0.0000 299.1500 0.6000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.2500 0.0000 298.3500 0.6000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.4500 0.0000 297.5500 0.6000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 296.6500 0.0000 296.7500 0.6000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.8500 0.0000 295.9500 0.6000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.0500 0.0000 295.1500 0.6000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 294.2500 0.0000 294.3500 0.6000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.4500 0.0000 293.5500 0.6000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.6500 0.0000 292.7500 0.6000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.8500 0.0000 291.9500 0.6000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.0500 0.0000 291.1500 0.6000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.2500 0.0000 290.3500 0.6000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.4500 0.0000 289.5500 0.6000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 288.6500 0.0000 288.7500 0.6000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.8500 0.0000 287.9500 0.6000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.0500 0.0000 287.1500 0.6000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.2500 0.0000 286.3500 0.6000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 285.4500 0.0000 285.5500 0.6000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 284.6500 0.0000 284.7500 0.6000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.8500 0.0000 283.9500 0.6000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.0500 0.0000 283.1500 0.6000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.2500 0.0000 282.3500 0.6000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.4500 0.0000 281.5500 0.6000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 280.6500 0.0000 280.7500 0.6000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.8500 0.0000 279.9500 0.6000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.0500 0.0000 279.1500 0.6000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 278.2500 0.0000 278.3500 0.6000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.4500 0.0000 277.5500 0.6000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.6500 0.0000 276.7500 0.6000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 275.8500 0.0000 275.9500 0.6000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 275.0500 0.0000 275.1500 0.6000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.2500 0.0000 274.3500 0.6000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 273.4500 0.0000 273.5500 0.6000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 272.6500 0.0000 272.7500 0.6000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.8500 0.0000 271.9500 0.6000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.0500 0.0000 271.1500 0.6000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 270.2500 0.0000 270.3500 0.6000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 269.4500 0.0000 269.5500 0.6000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 268.6500 0.0000 268.7500 0.6000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 267.8500 0.0000 267.9500 0.6000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 267.0500 0.0000 267.1500 0.6000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 266.2500 0.0000 266.3500 0.6000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 265.4500 0.0000 265.5500 0.6000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 264.6500 0.0000 264.7500 0.6000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 263.8500 0.0000 263.9500 0.6000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 263.0500 0.0000 263.1500 0.6000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 262.2500 0.0000 262.3500 0.6000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 261.4500 0.0000 261.5500 0.6000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 260.6500 0.0000 260.7500 0.6000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 259.8500 0.0000 259.9500 0.6000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 259.0500 0.0000 259.1500 0.6000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 258.2500 0.0000 258.3500 0.6000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 257.4500 0.0000 257.5500 0.6000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 256.6500 0.0000 256.7500 0.6000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.8500 0.0000 255.9500 0.6000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.0500 0.0000 255.1500 0.6000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 254.2500 0.0000 254.3500 0.6000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 253.4500 0.0000 253.5500 0.6000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.6500 0.0000 252.7500 0.6000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 251.8500 0.0000 251.9500 0.6000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 251.0500 0.0000 251.1500 0.6000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.2500 0.0000 250.3500 0.6000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 249.4500 0.0000 249.5500 0.6000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 248.6500 0.0000 248.7500 0.6000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.8500 0.0000 247.9500 0.6000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.0500 0.0000 247.1500 0.6000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 246.2500 0.0000 246.3500 0.6000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.4500 0.0000 245.5500 0.6000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.6500 0.0000 244.7500 0.6000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 243.8500 0.0000 243.9500 0.6000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 243.0500 0.0000 243.1500 0.6000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.2500 0.0000 242.3500 0.6000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 241.4500 0.0000 241.5500 0.6000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 240.6500 0.0000 240.7500 0.6000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.8500 0.0000 239.9500 0.6000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.0500 0.0000 239.1500 0.6000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 238.2500 0.0000 238.3500 0.6000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 237.4500 0.0000 237.5500 0.6000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.6500 0.0000 236.7500 0.6000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 235.8500 0.0000 235.9500 0.6000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 235.0500 0.0000 235.1500 0.6000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 234.2500 0.0000 234.3500 0.6000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.4500 0.0000 233.5500 0.6000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 232.6500 0.0000 232.7500 0.6000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.8500 0.0000 231.9500 0.6000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.0500 0.0000 231.1500 0.6000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 230.2500 0.0000 230.3500 0.6000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 229.4500 0.0000 229.5500 0.6000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.6500 0.0000 228.7500 0.6000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 227.8500 0.0000 227.9500 0.6000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 227.0500 0.0000 227.1500 0.6000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.2500 0.0000 226.3500 0.6000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.4500 0.0000 225.5500 0.6000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 224.6500 0.0000 224.7500 0.6000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.8500 0.0000 223.9500 0.6000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.0500 0.0000 223.1500 0.6000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 222.2500 0.0000 222.3500 0.6000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.4500 0.0000 221.5500 0.6000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.6500 0.0000 220.7500 0.6000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 219.8500 0.0000 219.9500 0.6000 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 199.7500 0.6000 199.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.9500 0.6000 199.0500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.1500 0.6000 198.2500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 197.3500 0.6000 197.4500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 196.5500 0.6000 196.6500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.7500 0.6000 195.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 194.9500 0.6000 195.0500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 194.1500 0.6000 194.2500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 193.3500 0.6000 193.4500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 192.5500 0.6000 192.6500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 191.7500 0.6000 191.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 190.9500 0.6000 191.0500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 190.1500 0.6000 190.2500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 189.3500 0.6000 189.4500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 188.5500 0.6000 188.6500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 187.7500 0.6000 187.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.9500 0.6000 187.0500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.1500 0.6000 186.2500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
    LAYER M3 ;
      RECT 0.0000 251.9500 438.8000 437.6000 ;
      RECT 0.7000 251.6500 438.8000 251.9500 ;
      RECT 0.0000 251.1500 438.8000 251.6500 ;
      RECT 0.7000 250.8500 438.8000 251.1500 ;
      RECT 0.0000 250.3500 438.8000 250.8500 ;
      RECT 0.7000 250.0500 438.8000 250.3500 ;
      RECT 0.0000 249.5500 438.8000 250.0500 ;
      RECT 0.7000 249.2500 438.8000 249.5500 ;
      RECT 0.0000 248.7500 438.8000 249.2500 ;
      RECT 0.7000 248.4500 438.8000 248.7500 ;
      RECT 0.0000 247.9500 438.8000 248.4500 ;
      RECT 0.7000 247.6500 438.8000 247.9500 ;
      RECT 0.0000 247.1500 438.8000 247.6500 ;
      RECT 0.7000 246.8500 438.8000 247.1500 ;
      RECT 0.0000 246.3500 438.8000 246.8500 ;
      RECT 0.7000 246.0500 438.8000 246.3500 ;
      RECT 0.0000 245.5500 438.8000 246.0500 ;
      RECT 0.7000 245.2500 438.8000 245.5500 ;
      RECT 0.0000 244.7500 438.8000 245.2500 ;
      RECT 0.7000 244.4500 438.8000 244.7500 ;
      RECT 0.0000 243.9500 438.8000 244.4500 ;
      RECT 0.7000 243.6500 438.8000 243.9500 ;
      RECT 0.0000 243.1500 438.8000 243.6500 ;
      RECT 0.7000 242.8500 438.8000 243.1500 ;
      RECT 0.0000 242.3500 438.8000 242.8500 ;
      RECT 0.7000 242.0500 438.8000 242.3500 ;
      RECT 0.0000 241.5500 438.8000 242.0500 ;
      RECT 0.7000 241.2500 438.8000 241.5500 ;
      RECT 0.0000 240.7500 438.8000 241.2500 ;
      RECT 0.7000 240.4500 438.8000 240.7500 ;
      RECT 0.0000 239.9500 438.8000 240.4500 ;
      RECT 0.7000 239.6500 438.8000 239.9500 ;
      RECT 0.0000 239.1500 438.8000 239.6500 ;
      RECT 0.7000 238.8500 438.8000 239.1500 ;
      RECT 0.0000 238.3500 438.8000 238.8500 ;
      RECT 0.7000 238.0500 438.8000 238.3500 ;
      RECT 0.0000 237.5500 438.8000 238.0500 ;
      RECT 0.7000 237.2500 438.8000 237.5500 ;
      RECT 0.0000 236.7500 438.8000 237.2500 ;
      RECT 0.7000 236.4500 438.8000 236.7500 ;
      RECT 0.0000 235.9500 438.8000 236.4500 ;
      RECT 0.7000 235.6500 438.8000 235.9500 ;
      RECT 0.0000 235.1500 438.8000 235.6500 ;
      RECT 0.7000 234.8500 438.8000 235.1500 ;
      RECT 0.0000 234.3500 438.8000 234.8500 ;
      RECT 0.7000 234.0500 438.8000 234.3500 ;
      RECT 0.0000 233.5500 438.8000 234.0500 ;
      RECT 0.7000 233.2500 438.8000 233.5500 ;
      RECT 0.0000 232.7500 438.8000 233.2500 ;
      RECT 0.7000 232.4500 438.8000 232.7500 ;
      RECT 0.0000 231.9500 438.8000 232.4500 ;
      RECT 0.7000 231.6500 438.8000 231.9500 ;
      RECT 0.0000 231.1500 438.8000 231.6500 ;
      RECT 0.7000 230.8500 438.8000 231.1500 ;
      RECT 0.0000 230.3500 438.8000 230.8500 ;
      RECT 0.7000 230.0500 438.8000 230.3500 ;
      RECT 0.0000 229.5500 438.8000 230.0500 ;
      RECT 0.7000 229.2500 438.8000 229.5500 ;
      RECT 0.0000 228.7500 438.8000 229.2500 ;
      RECT 0.7000 228.4500 438.8000 228.7500 ;
      RECT 0.0000 227.9500 438.8000 228.4500 ;
      RECT 0.7000 227.6500 438.8000 227.9500 ;
      RECT 0.0000 227.1500 438.8000 227.6500 ;
      RECT 0.7000 226.8500 438.8000 227.1500 ;
      RECT 0.0000 226.3500 438.8000 226.8500 ;
      RECT 0.7000 226.0500 438.8000 226.3500 ;
      RECT 0.0000 225.5500 438.8000 226.0500 ;
      RECT 0.7000 225.2500 438.8000 225.5500 ;
      RECT 0.0000 224.7500 438.8000 225.2500 ;
      RECT 0.7000 224.4500 438.8000 224.7500 ;
      RECT 0.0000 223.9500 438.8000 224.4500 ;
      RECT 0.7000 223.6500 438.8000 223.9500 ;
      RECT 0.0000 223.1500 438.8000 223.6500 ;
      RECT 0.7000 222.8500 438.8000 223.1500 ;
      RECT 0.0000 222.3500 438.8000 222.8500 ;
      RECT 0.7000 222.0500 438.8000 222.3500 ;
      RECT 0.0000 221.5500 438.8000 222.0500 ;
      RECT 0.7000 221.2500 438.8000 221.5500 ;
      RECT 0.0000 220.7500 438.8000 221.2500 ;
      RECT 0.7000 220.4500 438.8000 220.7500 ;
      RECT 0.0000 219.9500 438.8000 220.4500 ;
      RECT 0.7000 219.6500 438.8000 219.9500 ;
      RECT 0.0000 219.1500 438.8000 219.6500 ;
      RECT 0.7000 218.8500 438.8000 219.1500 ;
      RECT 0.0000 218.3500 438.8000 218.8500 ;
      RECT 0.7000 218.0500 438.8000 218.3500 ;
      RECT 0.0000 217.5500 438.8000 218.0500 ;
      RECT 0.7000 217.2500 438.8000 217.5500 ;
      RECT 0.0000 216.7500 438.8000 217.2500 ;
      RECT 0.7000 216.4500 438.8000 216.7500 ;
      RECT 0.0000 215.9500 438.8000 216.4500 ;
      RECT 0.7000 215.6500 438.8000 215.9500 ;
      RECT 0.0000 215.1500 438.8000 215.6500 ;
      RECT 0.7000 214.8500 438.8000 215.1500 ;
      RECT 0.0000 214.3500 438.8000 214.8500 ;
      RECT 0.7000 214.0500 438.8000 214.3500 ;
      RECT 0.0000 213.5500 438.8000 214.0500 ;
      RECT 0.7000 213.2500 438.8000 213.5500 ;
      RECT 0.0000 212.7500 438.8000 213.2500 ;
      RECT 0.7000 212.4500 438.8000 212.7500 ;
      RECT 0.0000 211.9500 438.8000 212.4500 ;
      RECT 0.7000 211.6500 438.8000 211.9500 ;
      RECT 0.0000 211.1500 438.8000 211.6500 ;
      RECT 0.7000 210.8500 438.8000 211.1500 ;
      RECT 0.0000 210.3500 438.8000 210.8500 ;
      RECT 0.7000 210.0500 438.8000 210.3500 ;
      RECT 0.0000 209.5500 438.8000 210.0500 ;
      RECT 0.7000 209.2500 438.8000 209.5500 ;
      RECT 0.0000 208.7500 438.8000 209.2500 ;
      RECT 0.7000 208.4500 438.8000 208.7500 ;
      RECT 0.0000 207.9500 438.8000 208.4500 ;
      RECT 0.7000 207.6500 438.8000 207.9500 ;
      RECT 0.0000 207.1500 438.8000 207.6500 ;
      RECT 0.7000 206.8500 438.8000 207.1500 ;
      RECT 0.0000 206.3500 438.8000 206.8500 ;
      RECT 0.7000 206.0500 438.8000 206.3500 ;
      RECT 0.0000 205.5500 438.8000 206.0500 ;
      RECT 0.7000 205.2500 438.8000 205.5500 ;
      RECT 0.0000 204.7500 438.8000 205.2500 ;
      RECT 0.7000 204.4500 438.8000 204.7500 ;
      RECT 0.0000 203.9500 438.8000 204.4500 ;
      RECT 0.7000 203.6500 438.8000 203.9500 ;
      RECT 0.0000 203.1500 438.8000 203.6500 ;
      RECT 0.7000 202.8500 438.8000 203.1500 ;
      RECT 0.0000 202.3500 438.8000 202.8500 ;
      RECT 0.7000 202.0500 438.8000 202.3500 ;
      RECT 0.0000 201.5500 438.8000 202.0500 ;
      RECT 0.7000 201.2500 438.8000 201.5500 ;
      RECT 0.0000 200.7500 438.8000 201.2500 ;
      RECT 0.7000 200.4500 438.8000 200.7500 ;
      RECT 0.0000 199.9500 438.8000 200.4500 ;
      RECT 0.7000 199.6500 438.8000 199.9500 ;
      RECT 0.0000 199.1500 438.8000 199.6500 ;
      RECT 0.7000 198.8500 438.8000 199.1500 ;
      RECT 0.0000 198.3500 438.8000 198.8500 ;
      RECT 0.7000 198.0500 438.8000 198.3500 ;
      RECT 0.0000 197.5500 438.8000 198.0500 ;
      RECT 0.7000 197.2500 438.8000 197.5500 ;
      RECT 0.0000 196.7500 438.8000 197.2500 ;
      RECT 0.7000 196.4500 438.8000 196.7500 ;
      RECT 0.0000 195.9500 438.8000 196.4500 ;
      RECT 0.7000 195.6500 438.8000 195.9500 ;
      RECT 0.0000 195.1500 438.8000 195.6500 ;
      RECT 0.7000 194.8500 438.8000 195.1500 ;
      RECT 0.0000 194.3500 438.8000 194.8500 ;
      RECT 0.7000 194.0500 438.8000 194.3500 ;
      RECT 0.0000 193.5500 438.8000 194.0500 ;
      RECT 0.7000 193.2500 438.8000 193.5500 ;
      RECT 0.0000 192.7500 438.8000 193.2500 ;
      RECT 0.7000 192.4500 438.8000 192.7500 ;
      RECT 0.0000 191.9500 438.8000 192.4500 ;
      RECT 0.7000 191.6500 438.8000 191.9500 ;
      RECT 0.0000 191.1500 438.8000 191.6500 ;
      RECT 0.7000 190.8500 438.8000 191.1500 ;
      RECT 0.0000 190.3500 438.8000 190.8500 ;
      RECT 0.7000 190.0500 438.8000 190.3500 ;
      RECT 0.0000 189.5500 438.8000 190.0500 ;
      RECT 0.7000 189.2500 438.8000 189.5500 ;
      RECT 0.0000 188.7500 438.8000 189.2500 ;
      RECT 0.7000 188.4500 438.8000 188.7500 ;
      RECT 0.0000 187.9500 438.8000 188.4500 ;
      RECT 0.7000 187.6500 438.8000 187.9500 ;
      RECT 0.0000 187.1500 438.8000 187.6500 ;
      RECT 0.7000 186.8500 438.8000 187.1500 ;
      RECT 0.0000 186.3500 438.8000 186.8500 ;
      RECT 0.7000 186.0500 438.8000 186.3500 ;
      RECT 0.0000 0.7600 438.8000 186.0500 ;
      RECT 347.3100 0.0000 438.8000 0.7600 ;
      RECT 346.5100 0.0000 346.8900 0.7600 ;
      RECT 345.7100 0.0000 346.0900 0.7600 ;
      RECT 344.9100 0.0000 345.2900 0.7600 ;
      RECT 344.1100 0.0000 344.4900 0.7600 ;
      RECT 343.3100 0.0000 343.6900 0.7600 ;
      RECT 342.5100 0.0000 342.8900 0.7600 ;
      RECT 341.7100 0.0000 342.0900 0.7600 ;
      RECT 340.9100 0.0000 341.2900 0.7600 ;
      RECT 340.1100 0.0000 340.4900 0.7600 ;
      RECT 339.3100 0.0000 339.6900 0.7600 ;
      RECT 338.5100 0.0000 338.8900 0.7600 ;
      RECT 337.7100 0.0000 338.0900 0.7600 ;
      RECT 336.9100 0.0000 337.2900 0.7600 ;
      RECT 336.1100 0.0000 336.4900 0.7600 ;
      RECT 335.3100 0.0000 335.6900 0.7600 ;
      RECT 334.5100 0.0000 334.8900 0.7600 ;
      RECT 333.7100 0.0000 334.0900 0.7600 ;
      RECT 332.9100 0.0000 333.2900 0.7600 ;
      RECT 332.1100 0.0000 332.4900 0.7600 ;
      RECT 331.3100 0.0000 331.6900 0.7600 ;
      RECT 330.5100 0.0000 330.8900 0.7600 ;
      RECT 329.7100 0.0000 330.0900 0.7600 ;
      RECT 328.9100 0.0000 329.2900 0.7600 ;
      RECT 328.1100 0.0000 328.4900 0.7600 ;
      RECT 327.3100 0.0000 327.6900 0.7600 ;
      RECT 326.5100 0.0000 326.8900 0.7600 ;
      RECT 325.7100 0.0000 326.0900 0.7600 ;
      RECT 324.9100 0.0000 325.2900 0.7600 ;
      RECT 324.1100 0.0000 324.4900 0.7600 ;
      RECT 323.3100 0.0000 323.6900 0.7600 ;
      RECT 322.5100 0.0000 322.8900 0.7600 ;
      RECT 321.7100 0.0000 322.0900 0.7600 ;
      RECT 320.9100 0.0000 321.2900 0.7600 ;
      RECT 320.1100 0.0000 320.4900 0.7600 ;
      RECT 319.3100 0.0000 319.6900 0.7600 ;
      RECT 318.5100 0.0000 318.8900 0.7600 ;
      RECT 317.7100 0.0000 318.0900 0.7600 ;
      RECT 316.9100 0.0000 317.2900 0.7600 ;
      RECT 316.1100 0.0000 316.4900 0.7600 ;
      RECT 315.3100 0.0000 315.6900 0.7600 ;
      RECT 314.5100 0.0000 314.8900 0.7600 ;
      RECT 313.7100 0.0000 314.0900 0.7600 ;
      RECT 312.9100 0.0000 313.2900 0.7600 ;
      RECT 312.1100 0.0000 312.4900 0.7600 ;
      RECT 311.3100 0.0000 311.6900 0.7600 ;
      RECT 310.5100 0.0000 310.8900 0.7600 ;
      RECT 309.7100 0.0000 310.0900 0.7600 ;
      RECT 308.9100 0.0000 309.2900 0.7600 ;
      RECT 308.1100 0.0000 308.4900 0.7600 ;
      RECT 307.3100 0.0000 307.6900 0.7600 ;
      RECT 306.5100 0.0000 306.8900 0.7600 ;
      RECT 305.7100 0.0000 306.0900 0.7600 ;
      RECT 304.9100 0.0000 305.2900 0.7600 ;
      RECT 304.1100 0.0000 304.4900 0.7600 ;
      RECT 303.3100 0.0000 303.6900 0.7600 ;
      RECT 302.5100 0.0000 302.8900 0.7600 ;
      RECT 301.7100 0.0000 302.0900 0.7600 ;
      RECT 300.9100 0.0000 301.2900 0.7600 ;
      RECT 300.1100 0.0000 300.4900 0.7600 ;
      RECT 299.3100 0.0000 299.6900 0.7600 ;
      RECT 298.5100 0.0000 298.8900 0.7600 ;
      RECT 297.7100 0.0000 298.0900 0.7600 ;
      RECT 296.9100 0.0000 297.2900 0.7600 ;
      RECT 296.1100 0.0000 296.4900 0.7600 ;
      RECT 295.3100 0.0000 295.6900 0.7600 ;
      RECT 294.5100 0.0000 294.8900 0.7600 ;
      RECT 293.7100 0.0000 294.0900 0.7600 ;
      RECT 292.9100 0.0000 293.2900 0.7600 ;
      RECT 292.1100 0.0000 292.4900 0.7600 ;
      RECT 291.3100 0.0000 291.6900 0.7600 ;
      RECT 290.5100 0.0000 290.8900 0.7600 ;
      RECT 289.7100 0.0000 290.0900 0.7600 ;
      RECT 288.9100 0.0000 289.2900 0.7600 ;
      RECT 288.1100 0.0000 288.4900 0.7600 ;
      RECT 287.3100 0.0000 287.6900 0.7600 ;
      RECT 286.5100 0.0000 286.8900 0.7600 ;
      RECT 285.7100 0.0000 286.0900 0.7600 ;
      RECT 284.9100 0.0000 285.2900 0.7600 ;
      RECT 284.1100 0.0000 284.4900 0.7600 ;
      RECT 283.3100 0.0000 283.6900 0.7600 ;
      RECT 282.5100 0.0000 282.8900 0.7600 ;
      RECT 281.7100 0.0000 282.0900 0.7600 ;
      RECT 280.9100 0.0000 281.2900 0.7600 ;
      RECT 280.1100 0.0000 280.4900 0.7600 ;
      RECT 279.3100 0.0000 279.6900 0.7600 ;
      RECT 278.5100 0.0000 278.8900 0.7600 ;
      RECT 277.7100 0.0000 278.0900 0.7600 ;
      RECT 276.9100 0.0000 277.2900 0.7600 ;
      RECT 276.1100 0.0000 276.4900 0.7600 ;
      RECT 275.3100 0.0000 275.6900 0.7600 ;
      RECT 274.5100 0.0000 274.8900 0.7600 ;
      RECT 273.7100 0.0000 274.0900 0.7600 ;
      RECT 272.9100 0.0000 273.2900 0.7600 ;
      RECT 272.1100 0.0000 272.4900 0.7600 ;
      RECT 271.3100 0.0000 271.6900 0.7600 ;
      RECT 270.5100 0.0000 270.8900 0.7600 ;
      RECT 269.7100 0.0000 270.0900 0.7600 ;
      RECT 268.9100 0.0000 269.2900 0.7600 ;
      RECT 268.1100 0.0000 268.4900 0.7600 ;
      RECT 267.3100 0.0000 267.6900 0.7600 ;
      RECT 266.5100 0.0000 266.8900 0.7600 ;
      RECT 265.7100 0.0000 266.0900 0.7600 ;
      RECT 264.9100 0.0000 265.2900 0.7600 ;
      RECT 264.1100 0.0000 264.4900 0.7600 ;
      RECT 263.3100 0.0000 263.6900 0.7600 ;
      RECT 262.5100 0.0000 262.8900 0.7600 ;
      RECT 261.7100 0.0000 262.0900 0.7600 ;
      RECT 260.9100 0.0000 261.2900 0.7600 ;
      RECT 260.1100 0.0000 260.4900 0.7600 ;
      RECT 259.3100 0.0000 259.6900 0.7600 ;
      RECT 258.5100 0.0000 258.8900 0.7600 ;
      RECT 257.7100 0.0000 258.0900 0.7600 ;
      RECT 256.9100 0.0000 257.2900 0.7600 ;
      RECT 256.1100 0.0000 256.4900 0.7600 ;
      RECT 255.3100 0.0000 255.6900 0.7600 ;
      RECT 254.5100 0.0000 254.8900 0.7600 ;
      RECT 253.7100 0.0000 254.0900 0.7600 ;
      RECT 252.9100 0.0000 253.2900 0.7600 ;
      RECT 252.1100 0.0000 252.4900 0.7600 ;
      RECT 251.3100 0.0000 251.6900 0.7600 ;
      RECT 250.5100 0.0000 250.8900 0.7600 ;
      RECT 249.7100 0.0000 250.0900 0.7600 ;
      RECT 248.9100 0.0000 249.2900 0.7600 ;
      RECT 248.1100 0.0000 248.4900 0.7600 ;
      RECT 247.3100 0.0000 247.6900 0.7600 ;
      RECT 246.5100 0.0000 246.8900 0.7600 ;
      RECT 245.7100 0.0000 246.0900 0.7600 ;
      RECT 244.9100 0.0000 245.2900 0.7600 ;
      RECT 244.1100 0.0000 244.4900 0.7600 ;
      RECT 243.3100 0.0000 243.6900 0.7600 ;
      RECT 242.5100 0.0000 242.8900 0.7600 ;
      RECT 241.7100 0.0000 242.0900 0.7600 ;
      RECT 240.9100 0.0000 241.2900 0.7600 ;
      RECT 240.1100 0.0000 240.4900 0.7600 ;
      RECT 239.3100 0.0000 239.6900 0.7600 ;
      RECT 238.5100 0.0000 238.8900 0.7600 ;
      RECT 237.7100 0.0000 238.0900 0.7600 ;
      RECT 236.9100 0.0000 237.2900 0.7600 ;
      RECT 236.1100 0.0000 236.4900 0.7600 ;
      RECT 235.3100 0.0000 235.6900 0.7600 ;
      RECT 234.5100 0.0000 234.8900 0.7600 ;
      RECT 233.7100 0.0000 234.0900 0.7600 ;
      RECT 232.9100 0.0000 233.2900 0.7600 ;
      RECT 232.1100 0.0000 232.4900 0.7600 ;
      RECT 231.3100 0.0000 231.6900 0.7600 ;
      RECT 230.5100 0.0000 230.8900 0.7600 ;
      RECT 229.7100 0.0000 230.0900 0.7600 ;
      RECT 228.9100 0.0000 229.2900 0.7600 ;
      RECT 228.1100 0.0000 228.4900 0.7600 ;
      RECT 227.3100 0.0000 227.6900 0.7600 ;
      RECT 226.5100 0.0000 226.8900 0.7600 ;
      RECT 225.7100 0.0000 226.0900 0.7600 ;
      RECT 224.9100 0.0000 225.2900 0.7600 ;
      RECT 224.1100 0.0000 224.4900 0.7600 ;
      RECT 223.3100 0.0000 223.6900 0.7600 ;
      RECT 222.5100 0.0000 222.8900 0.7600 ;
      RECT 221.7100 0.0000 222.0900 0.7600 ;
      RECT 220.9100 0.0000 221.2900 0.7600 ;
      RECT 220.1100 0.0000 220.4900 0.7600 ;
      RECT 219.3100 0.0000 219.6900 0.7600 ;
      RECT 218.5100 0.0000 218.8900 0.7600 ;
      RECT 217.7100 0.0000 218.0900 0.7600 ;
      RECT 216.9100 0.0000 217.2900 0.7600 ;
      RECT 216.1100 0.0000 216.4900 0.7600 ;
      RECT 215.3100 0.0000 215.6900 0.7600 ;
      RECT 214.5100 0.0000 214.8900 0.7600 ;
      RECT 213.7100 0.0000 214.0900 0.7600 ;
      RECT 212.9100 0.0000 213.2900 0.7600 ;
      RECT 212.1100 0.0000 212.4900 0.7600 ;
      RECT 211.3100 0.0000 211.6900 0.7600 ;
      RECT 210.5100 0.0000 210.8900 0.7600 ;
      RECT 209.7100 0.0000 210.0900 0.7600 ;
      RECT 208.9100 0.0000 209.2900 0.7600 ;
      RECT 208.1100 0.0000 208.4900 0.7600 ;
      RECT 207.3100 0.0000 207.6900 0.7600 ;
      RECT 206.5100 0.0000 206.8900 0.7600 ;
      RECT 205.7100 0.0000 206.0900 0.7600 ;
      RECT 204.9100 0.0000 205.2900 0.7600 ;
      RECT 204.1100 0.0000 204.4900 0.7600 ;
      RECT 203.3100 0.0000 203.6900 0.7600 ;
      RECT 202.5100 0.0000 202.8900 0.7600 ;
      RECT 201.7100 0.0000 202.0900 0.7600 ;
      RECT 200.9100 0.0000 201.2900 0.7600 ;
      RECT 200.1100 0.0000 200.4900 0.7600 ;
      RECT 199.3100 0.0000 199.6900 0.7600 ;
      RECT 198.5100 0.0000 198.8900 0.7600 ;
      RECT 197.7100 0.0000 198.0900 0.7600 ;
      RECT 196.9100 0.0000 197.2900 0.7600 ;
      RECT 196.1100 0.0000 196.4900 0.7600 ;
      RECT 195.3100 0.0000 195.6900 0.7600 ;
      RECT 194.5100 0.0000 194.8900 0.7600 ;
      RECT 193.7100 0.0000 194.0900 0.7600 ;
      RECT 192.9100 0.0000 193.2900 0.7600 ;
      RECT 192.1100 0.0000 192.4900 0.7600 ;
      RECT 191.3100 0.0000 191.6900 0.7600 ;
      RECT 190.5100 0.0000 190.8900 0.7600 ;
      RECT 189.7100 0.0000 190.0900 0.7600 ;
      RECT 188.9100 0.0000 189.2900 0.7600 ;
      RECT 188.1100 0.0000 188.4900 0.7600 ;
      RECT 187.3100 0.0000 187.6900 0.7600 ;
      RECT 186.5100 0.0000 186.8900 0.7600 ;
      RECT 185.7100 0.0000 186.0900 0.7600 ;
      RECT 184.9100 0.0000 185.2900 0.7600 ;
      RECT 184.1100 0.0000 184.4900 0.7600 ;
      RECT 183.3100 0.0000 183.6900 0.7600 ;
      RECT 182.5100 0.0000 182.8900 0.7600 ;
      RECT 181.7100 0.0000 182.0900 0.7600 ;
      RECT 180.9100 0.0000 181.2900 0.7600 ;
      RECT 180.1100 0.0000 180.4900 0.7600 ;
      RECT 179.3100 0.0000 179.6900 0.7600 ;
      RECT 178.5100 0.0000 178.8900 0.7600 ;
      RECT 177.7100 0.0000 178.0900 0.7600 ;
      RECT 176.9100 0.0000 177.2900 0.7600 ;
      RECT 176.1100 0.0000 176.4900 0.7600 ;
      RECT 175.3100 0.0000 175.6900 0.7600 ;
      RECT 174.5100 0.0000 174.8900 0.7600 ;
      RECT 173.7100 0.0000 174.0900 0.7600 ;
      RECT 172.9100 0.0000 173.2900 0.7600 ;
      RECT 172.1100 0.0000 172.4900 0.7600 ;
      RECT 171.3100 0.0000 171.6900 0.7600 ;
      RECT 170.5100 0.0000 170.8900 0.7600 ;
      RECT 169.7100 0.0000 170.0900 0.7600 ;
      RECT 168.9100 0.0000 169.2900 0.7600 ;
      RECT 168.1100 0.0000 168.4900 0.7600 ;
      RECT 167.3100 0.0000 167.6900 0.7600 ;
      RECT 166.5100 0.0000 166.8900 0.7600 ;
      RECT 165.7100 0.0000 166.0900 0.7600 ;
      RECT 164.9100 0.0000 165.2900 0.7600 ;
      RECT 164.1100 0.0000 164.4900 0.7600 ;
      RECT 163.3100 0.0000 163.6900 0.7600 ;
      RECT 162.5100 0.0000 162.8900 0.7600 ;
      RECT 161.7100 0.0000 162.0900 0.7600 ;
      RECT 160.9100 0.0000 161.2900 0.7600 ;
      RECT 160.1100 0.0000 160.4900 0.7600 ;
      RECT 159.3100 0.0000 159.6900 0.7600 ;
      RECT 158.5100 0.0000 158.8900 0.7600 ;
      RECT 157.7100 0.0000 158.0900 0.7600 ;
      RECT 156.9100 0.0000 157.2900 0.7600 ;
      RECT 156.1100 0.0000 156.4900 0.7600 ;
      RECT 155.3100 0.0000 155.6900 0.7600 ;
      RECT 154.5100 0.0000 154.8900 0.7600 ;
      RECT 153.7100 0.0000 154.0900 0.7600 ;
      RECT 152.9100 0.0000 153.2900 0.7600 ;
      RECT 152.1100 0.0000 152.4900 0.7600 ;
      RECT 151.3100 0.0000 151.6900 0.7600 ;
      RECT 150.5100 0.0000 150.8900 0.7600 ;
      RECT 149.7100 0.0000 150.0900 0.7600 ;
      RECT 148.9100 0.0000 149.2900 0.7600 ;
      RECT 148.1100 0.0000 148.4900 0.7600 ;
      RECT 147.3100 0.0000 147.6900 0.7600 ;
      RECT 146.5100 0.0000 146.8900 0.7600 ;
      RECT 145.7100 0.0000 146.0900 0.7600 ;
      RECT 144.9100 0.0000 145.2900 0.7600 ;
      RECT 144.1100 0.0000 144.4900 0.7600 ;
      RECT 143.3100 0.0000 143.6900 0.7600 ;
      RECT 142.5100 0.0000 142.8900 0.7600 ;
      RECT 141.7100 0.0000 142.0900 0.7600 ;
      RECT 140.9100 0.0000 141.2900 0.7600 ;
      RECT 140.1100 0.0000 140.4900 0.7600 ;
      RECT 139.3100 0.0000 139.6900 0.7600 ;
      RECT 138.5100 0.0000 138.8900 0.7600 ;
      RECT 137.7100 0.0000 138.0900 0.7600 ;
      RECT 136.9100 0.0000 137.2900 0.7600 ;
      RECT 136.1100 0.0000 136.4900 0.7600 ;
      RECT 135.3100 0.0000 135.6900 0.7600 ;
      RECT 134.5100 0.0000 134.8900 0.7600 ;
      RECT 133.7100 0.0000 134.0900 0.7600 ;
      RECT 132.9100 0.0000 133.2900 0.7600 ;
      RECT 132.1100 0.0000 132.4900 0.7600 ;
      RECT 131.3100 0.0000 131.6900 0.7600 ;
      RECT 130.5100 0.0000 130.8900 0.7600 ;
      RECT 129.7100 0.0000 130.0900 0.7600 ;
      RECT 128.9100 0.0000 129.2900 0.7600 ;
      RECT 128.1100 0.0000 128.4900 0.7600 ;
      RECT 127.3100 0.0000 127.6900 0.7600 ;
      RECT 126.5100 0.0000 126.8900 0.7600 ;
      RECT 125.7100 0.0000 126.0900 0.7600 ;
      RECT 124.9100 0.0000 125.2900 0.7600 ;
      RECT 124.1100 0.0000 124.4900 0.7600 ;
      RECT 123.3100 0.0000 123.6900 0.7600 ;
      RECT 122.5100 0.0000 122.8900 0.7600 ;
      RECT 121.7100 0.0000 122.0900 0.7600 ;
      RECT 120.9100 0.0000 121.2900 0.7600 ;
      RECT 120.1100 0.0000 120.4900 0.7600 ;
      RECT 119.3100 0.0000 119.6900 0.7600 ;
      RECT 118.5100 0.0000 118.8900 0.7600 ;
      RECT 117.7100 0.0000 118.0900 0.7600 ;
      RECT 116.9100 0.0000 117.2900 0.7600 ;
      RECT 116.1100 0.0000 116.4900 0.7600 ;
      RECT 115.3100 0.0000 115.6900 0.7600 ;
      RECT 114.5100 0.0000 114.8900 0.7600 ;
      RECT 113.7100 0.0000 114.0900 0.7600 ;
      RECT 112.9100 0.0000 113.2900 0.7600 ;
      RECT 112.1100 0.0000 112.4900 0.7600 ;
      RECT 111.3100 0.0000 111.6900 0.7600 ;
      RECT 110.5100 0.0000 110.8900 0.7600 ;
      RECT 109.7100 0.0000 110.0900 0.7600 ;
      RECT 108.9100 0.0000 109.2900 0.7600 ;
      RECT 108.1100 0.0000 108.4900 0.7600 ;
      RECT 107.3100 0.0000 107.6900 0.7600 ;
      RECT 106.5100 0.0000 106.8900 0.7600 ;
      RECT 105.7100 0.0000 106.0900 0.7600 ;
      RECT 104.9100 0.0000 105.2900 0.7600 ;
      RECT 104.1100 0.0000 104.4900 0.7600 ;
      RECT 103.3100 0.0000 103.6900 0.7600 ;
      RECT 102.5100 0.0000 102.8900 0.7600 ;
      RECT 101.7100 0.0000 102.0900 0.7600 ;
      RECT 100.9100 0.0000 101.2900 0.7600 ;
      RECT 100.1100 0.0000 100.4900 0.7600 ;
      RECT 99.3100 0.0000 99.6900 0.7600 ;
      RECT 98.5100 0.0000 98.8900 0.7600 ;
      RECT 97.7100 0.0000 98.0900 0.7600 ;
      RECT 96.9100 0.0000 97.2900 0.7600 ;
      RECT 96.1100 0.0000 96.4900 0.7600 ;
      RECT 95.3100 0.0000 95.6900 0.7600 ;
      RECT 94.5100 0.0000 94.8900 0.7600 ;
      RECT 93.7100 0.0000 94.0900 0.7600 ;
      RECT 92.9100 0.0000 93.2900 0.7600 ;
      RECT 92.1100 0.0000 92.4900 0.7600 ;
      RECT 0.0000 0.0000 91.6900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 438.8000 437.6000 ;
  END
END core

END LIBRARY
