##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 08:13:47 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 118.4000 BY 115.4000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.5500 0.6000 45.6500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.0500 0.0000 10.1500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.8500 0.0000 10.9500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.6500 0.0000 11.7500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.4500 0.0000 12.5500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.2500 0.0000 13.3500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.0500 0.0000 14.1500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.8500 0.0000 14.9500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6500 0.0000 15.7500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4500 0.0000 16.5500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.2500 0.0000 17.3500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.0500 0.0000 18.1500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.8500 0.0000 18.9500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.6500 0.0000 19.7500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4500 0.0000 20.5500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.2500 0.0000 21.3500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.0500 0.0000 22.1500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.8500 0.0000 22.9500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.6500 0.0000 23.7500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.4500 0.0000 24.5500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2500 0.0000 25.3500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.0500 0.0000 26.1500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.8500 0.0000 26.9500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.6500 0.0000 27.7500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4500 0.0000 28.5500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2500 0.0000 29.3500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.0500 0.0000 30.1500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.8500 0.0000 30.9500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.6500 0.0000 31.7500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4500 0.0000 32.5500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.2500 0.0000 33.3500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.0500 0.0000 34.1500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.8500 0.0000 34.9500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.6500 0.0000 35.7500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.4500 0.0000 36.5500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.2500 0.0000 37.3500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0500 0.0000 38.1500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.8500 0.0000 38.9500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.6500 0.0000 39.7500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.4500 0.0000 40.5500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.2500 0.0000 41.3500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.0500 0.0000 42.1500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.8500 0.0000 42.9500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.6500 0.0000 43.7500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.4500 0.0000 44.5500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.2500 0.0000 45.3500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.0500 0.0000 46.1500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8500 0.0000 46.9500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.6500 0.0000 47.7500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.4500 0.0000 48.5500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.2500 0.0000 49.3500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.0500 0.0000 50.1500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8500 0.0000 50.9500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.6500 0.0000 51.7500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.4500 0.0000 52.5500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.2500 0.0000 53.3500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.0500 0.0000 54.1500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.8500 0.0000 54.9500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.6500 0.0000 55.7500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.4500 0.0000 56.5500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.2500 0.0000 57.3500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.0500 0.0000 58.1500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8500 0.0000 58.9500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.6500 0.0000 59.7500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.4500 0.0000 60.5500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.2500 0.0000 61.3500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.0500 0.0000 62.1500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8500 0.0000 62.9500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.6500 0.0000 63.7500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.4500 0.0000 64.5500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.2500 0.0000 65.3500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.0500 0.0000 66.1500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 0.0000 66.9500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.6500 0.0000 67.7500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.4500 0.0000 68.5500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.2500 0.0000 69.3500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.0500 0.0000 70.1500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8500 0.0000 70.9500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.6500 0.0000 71.7500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.4500 0.0000 72.5500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.2500 0.0000 73.3500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 0.0000 74.1500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.8500 0.0000 74.9500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.6500 0.0000 75.7500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.4500 0.0000 76.5500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.2500 0.0000 77.3500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.0500 0.0000 78.1500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8500 0.0000 78.9500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.6500 0.0000 79.7500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.4500 0.0000 80.5500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.2500 0.0000 81.3500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.0500 0.0000 82.1500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.8500 0.0000 82.9500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.6500 0.0000 83.7500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.4500 0.0000 84.5500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.2500 0.0000 85.3500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.0500 0.0000 86.1500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.8500 0.0000 86.9500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.6500 0.0000 87.7500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.4500 0.0000 88.5500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.2500 0.0000 89.3500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.0500 0.0000 90.1500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 0.0000 90.9500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.6500 0.0000 91.7500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.4500 0.0000 92.5500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.2500 0.0000 93.3500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 0.0000 94.1500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 0.0000 94.9500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.6500 0.0000 95.7500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.4500 0.0000 96.5500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.2500 0.0000 97.3500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 0.0000 98.1500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 0.0000 98.9500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.6500 0.0000 99.7500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.4500 0.0000 100.5500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.2500 0.0000 101.3500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 0.0000 102.1500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 0.0000 102.9500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.6500 0.0000 103.7500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.4500 0.0000 104.5500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.2500 0.0000 105.3500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 0.0000 106.1500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 0.0000 106.9500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.6500 0.0000 107.7500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 0.0000 108.5500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.2500 0.0000 109.3500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 0.0000 110.1500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 0.0000 110.9500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.6500 0.0000 111.7500 0.6000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.0500 114.8000 10.1500 115.4000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.8500 114.8000 10.9500 115.4000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.6500 114.8000 11.7500 115.4000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.4500 114.8000 12.5500 115.4000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.2500 114.8000 13.3500 115.4000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.0500 114.8000 14.1500 115.4000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.8500 114.8000 14.9500 115.4000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.6500 114.8000 15.7500 115.4000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4500 114.8000 16.5500 115.4000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.2500 114.8000 17.3500 115.4000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.0500 114.8000 18.1500 115.4000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.8500 114.8000 18.9500 115.4000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.6500 114.8000 19.7500 115.4000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.4500 114.8000 20.5500 115.4000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.2500 114.8000 21.3500 115.4000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.0500 114.8000 22.1500 115.4000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.8500 114.8000 22.9500 115.4000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.6500 114.8000 23.7500 115.4000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.4500 114.8000 24.5500 115.4000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.2500 114.8000 25.3500 115.4000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.0500 114.8000 26.1500 115.4000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.8500 114.8000 26.9500 115.4000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.6500 114.8000 27.7500 115.4000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4500 114.8000 28.5500 115.4000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.2500 114.8000 29.3500 115.4000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.0500 114.8000 30.1500 115.4000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.8500 114.8000 30.9500 115.4000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.6500 114.8000 31.7500 115.4000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4500 114.8000 32.5500 115.4000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.2500 114.8000 33.3500 115.4000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.0500 114.8000 34.1500 115.4000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.8500 114.8000 34.9500 115.4000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.6500 114.8000 35.7500 115.4000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.4500 114.8000 36.5500 115.4000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.2500 114.8000 37.3500 115.4000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0500 114.8000 38.1500 115.4000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.8500 114.8000 38.9500 115.4000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.6500 114.8000 39.7500 115.4000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.4500 114.8000 40.5500 115.4000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.2500 114.8000 41.3500 115.4000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.0500 114.8000 42.1500 115.4000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.8500 114.8000 42.9500 115.4000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.6500 114.8000 43.7500 115.4000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.4500 114.8000 44.5500 115.4000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.2500 114.8000 45.3500 115.4000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.0500 114.8000 46.1500 115.4000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8500 114.8000 46.9500 115.4000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.6500 114.8000 47.7500 115.4000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.4500 114.8000 48.5500 115.4000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.2500 114.8000 49.3500 115.4000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.0500 114.8000 50.1500 115.4000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8500 114.8000 50.9500 115.4000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.6500 114.8000 51.7500 115.4000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.4500 114.8000 52.5500 115.4000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.2500 114.8000 53.3500 115.4000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.0500 114.8000 54.1500 115.4000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.8500 114.8000 54.9500 115.4000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.6500 114.8000 55.7500 115.4000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.4500 114.8000 56.5500 115.4000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.2500 114.8000 57.3500 115.4000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.0500 114.8000 58.1500 115.4000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8500 114.8000 58.9500 115.4000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.6500 114.8000 59.7500 115.4000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.4500 114.8000 60.5500 115.4000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.2500 114.8000 61.3500 115.4000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.0500 114.8000 62.1500 115.4000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8500 114.8000 62.9500 115.4000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.6500 114.8000 63.7500 115.4000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.4500 114.8000 64.5500 115.4000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.2500 114.8000 65.3500 115.4000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.0500 114.8000 66.1500 115.4000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 114.8000 66.9500 115.4000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.6500 114.8000 67.7500 115.4000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.4500 114.8000 68.5500 115.4000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.2500 114.8000 69.3500 115.4000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.0500 114.8000 70.1500 115.4000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8500 114.8000 70.9500 115.4000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.6500 114.8000 71.7500 115.4000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.4500 114.8000 72.5500 115.4000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.2500 114.8000 73.3500 115.4000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 114.8000 74.1500 115.4000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.8500 114.8000 74.9500 115.4000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.6500 114.8000 75.7500 115.4000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.4500 114.8000 76.5500 115.4000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.2500 114.8000 77.3500 115.4000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.0500 114.8000 78.1500 115.4000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8500 114.8000 78.9500 115.4000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.6500 114.8000 79.7500 115.4000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.4500 114.8000 80.5500 115.4000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.2500 114.8000 81.3500 115.4000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.0500 114.8000 82.1500 115.4000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.8500 114.8000 82.9500 115.4000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.6500 114.8000 83.7500 115.4000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.4500 114.8000 84.5500 115.4000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.2500 114.8000 85.3500 115.4000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.0500 114.8000 86.1500 115.4000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.8500 114.8000 86.9500 115.4000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.6500 114.8000 87.7500 115.4000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.4500 114.8000 88.5500 115.4000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.2500 114.8000 89.3500 115.4000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.0500 114.8000 90.1500 115.4000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 114.8000 90.9500 115.4000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.6500 114.8000 91.7500 115.4000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.4500 114.8000 92.5500 115.4000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.2500 114.8000 93.3500 115.4000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 114.8000 94.1500 115.4000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 114.8000 94.9500 115.4000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.6500 114.8000 95.7500 115.4000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.4500 114.8000 96.5500 115.4000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.2500 114.8000 97.3500 115.4000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 114.8000 98.1500 115.4000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 114.8000 98.9500 115.4000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.6500 114.8000 99.7500 115.4000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.4500 114.8000 100.5500 115.4000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.2500 114.8000 101.3500 115.4000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 114.8000 102.1500 115.4000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 114.8000 102.9500 115.4000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.6500 114.8000 103.7500 115.4000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.4500 114.8000 104.5500 115.4000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.2500 114.8000 105.3500 115.4000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 114.8000 106.1500 115.4000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 114.8000 106.9500 115.4000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.6500 114.8000 107.7500 115.4000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 114.8000 108.5500 115.4000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.2500 114.8000 109.3500 115.4000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 114.8000 110.1500 115.4000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 114.8000 110.9500 115.4000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.6500 114.8000 111.7500 115.4000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.5500 0.6000 65.6500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 69.5500 0.6000 69.6500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.5500 0.6000 49.6500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.5500 0.6000 53.6500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.5500 0.6000 57.6500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.5500 0.6000 61.6500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 7.0000 1.0000 8.0000 114.4000 ;
        RECT 114.0000 1.0000 115.0000 114.4000 ;
        RECT 7.0000 114.2350 8.0000 114.5650 ;
        RECT 114.0000 114.2350 115.0000 114.5650 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 5.0000 1.0000 6.0000 114.4000 ;
        RECT 112.0000 1.0000 113.0000 114.4000 ;
        RECT 5.0000 0.8350 6.0000 1.1650 ;
        RECT 112.0000 0.8350 113.0000 1.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 118.4000 115.4000 ;
    LAYER M2 ;
      RECT 111.8500 114.7000 118.4000 115.4000 ;
      RECT 111.0500 114.7000 111.5500 115.4000 ;
      RECT 110.2500 114.7000 110.7500 115.4000 ;
      RECT 109.4500 114.7000 109.9500 115.4000 ;
      RECT 108.6500 114.7000 109.1500 115.4000 ;
      RECT 107.8500 114.7000 108.3500 115.4000 ;
      RECT 107.0500 114.7000 107.5500 115.4000 ;
      RECT 106.2500 114.7000 106.7500 115.4000 ;
      RECT 105.4500 114.7000 105.9500 115.4000 ;
      RECT 104.6500 114.7000 105.1500 115.4000 ;
      RECT 103.8500 114.7000 104.3500 115.4000 ;
      RECT 103.0500 114.7000 103.5500 115.4000 ;
      RECT 102.2500 114.7000 102.7500 115.4000 ;
      RECT 101.4500 114.7000 101.9500 115.4000 ;
      RECT 100.6500 114.7000 101.1500 115.4000 ;
      RECT 99.8500 114.7000 100.3500 115.4000 ;
      RECT 99.0500 114.7000 99.5500 115.4000 ;
      RECT 98.2500 114.7000 98.7500 115.4000 ;
      RECT 97.4500 114.7000 97.9500 115.4000 ;
      RECT 96.6500 114.7000 97.1500 115.4000 ;
      RECT 95.8500 114.7000 96.3500 115.4000 ;
      RECT 95.0500 114.7000 95.5500 115.4000 ;
      RECT 94.2500 114.7000 94.7500 115.4000 ;
      RECT 93.4500 114.7000 93.9500 115.4000 ;
      RECT 92.6500 114.7000 93.1500 115.4000 ;
      RECT 91.8500 114.7000 92.3500 115.4000 ;
      RECT 91.0500 114.7000 91.5500 115.4000 ;
      RECT 90.2500 114.7000 90.7500 115.4000 ;
      RECT 89.4500 114.7000 89.9500 115.4000 ;
      RECT 88.6500 114.7000 89.1500 115.4000 ;
      RECT 87.8500 114.7000 88.3500 115.4000 ;
      RECT 87.0500 114.7000 87.5500 115.4000 ;
      RECT 86.2500 114.7000 86.7500 115.4000 ;
      RECT 85.4500 114.7000 85.9500 115.4000 ;
      RECT 84.6500 114.7000 85.1500 115.4000 ;
      RECT 83.8500 114.7000 84.3500 115.4000 ;
      RECT 83.0500 114.7000 83.5500 115.4000 ;
      RECT 82.2500 114.7000 82.7500 115.4000 ;
      RECT 81.4500 114.7000 81.9500 115.4000 ;
      RECT 80.6500 114.7000 81.1500 115.4000 ;
      RECT 79.8500 114.7000 80.3500 115.4000 ;
      RECT 79.0500 114.7000 79.5500 115.4000 ;
      RECT 78.2500 114.7000 78.7500 115.4000 ;
      RECT 77.4500 114.7000 77.9500 115.4000 ;
      RECT 76.6500 114.7000 77.1500 115.4000 ;
      RECT 75.8500 114.7000 76.3500 115.4000 ;
      RECT 75.0500 114.7000 75.5500 115.4000 ;
      RECT 74.2500 114.7000 74.7500 115.4000 ;
      RECT 73.4500 114.7000 73.9500 115.4000 ;
      RECT 72.6500 114.7000 73.1500 115.4000 ;
      RECT 71.8500 114.7000 72.3500 115.4000 ;
      RECT 71.0500 114.7000 71.5500 115.4000 ;
      RECT 70.2500 114.7000 70.7500 115.4000 ;
      RECT 69.4500 114.7000 69.9500 115.4000 ;
      RECT 68.6500 114.7000 69.1500 115.4000 ;
      RECT 67.8500 114.7000 68.3500 115.4000 ;
      RECT 67.0500 114.7000 67.5500 115.4000 ;
      RECT 66.2500 114.7000 66.7500 115.4000 ;
      RECT 65.4500 114.7000 65.9500 115.4000 ;
      RECT 64.6500 114.7000 65.1500 115.4000 ;
      RECT 63.8500 114.7000 64.3500 115.4000 ;
      RECT 63.0500 114.7000 63.5500 115.4000 ;
      RECT 62.2500 114.7000 62.7500 115.4000 ;
      RECT 61.4500 114.7000 61.9500 115.4000 ;
      RECT 60.6500 114.7000 61.1500 115.4000 ;
      RECT 59.8500 114.7000 60.3500 115.4000 ;
      RECT 59.0500 114.7000 59.5500 115.4000 ;
      RECT 58.2500 114.7000 58.7500 115.4000 ;
      RECT 57.4500 114.7000 57.9500 115.4000 ;
      RECT 56.6500 114.7000 57.1500 115.4000 ;
      RECT 55.8500 114.7000 56.3500 115.4000 ;
      RECT 55.0500 114.7000 55.5500 115.4000 ;
      RECT 54.2500 114.7000 54.7500 115.4000 ;
      RECT 53.4500 114.7000 53.9500 115.4000 ;
      RECT 52.6500 114.7000 53.1500 115.4000 ;
      RECT 51.8500 114.7000 52.3500 115.4000 ;
      RECT 51.0500 114.7000 51.5500 115.4000 ;
      RECT 50.2500 114.7000 50.7500 115.4000 ;
      RECT 49.4500 114.7000 49.9500 115.4000 ;
      RECT 48.6500 114.7000 49.1500 115.4000 ;
      RECT 47.8500 114.7000 48.3500 115.4000 ;
      RECT 47.0500 114.7000 47.5500 115.4000 ;
      RECT 46.2500 114.7000 46.7500 115.4000 ;
      RECT 45.4500 114.7000 45.9500 115.4000 ;
      RECT 44.6500 114.7000 45.1500 115.4000 ;
      RECT 43.8500 114.7000 44.3500 115.4000 ;
      RECT 43.0500 114.7000 43.5500 115.4000 ;
      RECT 42.2500 114.7000 42.7500 115.4000 ;
      RECT 41.4500 114.7000 41.9500 115.4000 ;
      RECT 40.6500 114.7000 41.1500 115.4000 ;
      RECT 39.8500 114.7000 40.3500 115.4000 ;
      RECT 39.0500 114.7000 39.5500 115.4000 ;
      RECT 38.2500 114.7000 38.7500 115.4000 ;
      RECT 37.4500 114.7000 37.9500 115.4000 ;
      RECT 36.6500 114.7000 37.1500 115.4000 ;
      RECT 35.8500 114.7000 36.3500 115.4000 ;
      RECT 35.0500 114.7000 35.5500 115.4000 ;
      RECT 34.2500 114.7000 34.7500 115.4000 ;
      RECT 33.4500 114.7000 33.9500 115.4000 ;
      RECT 32.6500 114.7000 33.1500 115.4000 ;
      RECT 31.8500 114.7000 32.3500 115.4000 ;
      RECT 31.0500 114.7000 31.5500 115.4000 ;
      RECT 30.2500 114.7000 30.7500 115.4000 ;
      RECT 29.4500 114.7000 29.9500 115.4000 ;
      RECT 28.6500 114.7000 29.1500 115.4000 ;
      RECT 27.8500 114.7000 28.3500 115.4000 ;
      RECT 27.0500 114.7000 27.5500 115.4000 ;
      RECT 26.2500 114.7000 26.7500 115.4000 ;
      RECT 25.4500 114.7000 25.9500 115.4000 ;
      RECT 24.6500 114.7000 25.1500 115.4000 ;
      RECT 23.8500 114.7000 24.3500 115.4000 ;
      RECT 23.0500 114.7000 23.5500 115.4000 ;
      RECT 22.2500 114.7000 22.7500 115.4000 ;
      RECT 21.4500 114.7000 21.9500 115.4000 ;
      RECT 20.6500 114.7000 21.1500 115.4000 ;
      RECT 19.8500 114.7000 20.3500 115.4000 ;
      RECT 19.0500 114.7000 19.5500 115.4000 ;
      RECT 18.2500 114.7000 18.7500 115.4000 ;
      RECT 17.4500 114.7000 17.9500 115.4000 ;
      RECT 16.6500 114.7000 17.1500 115.4000 ;
      RECT 15.8500 114.7000 16.3500 115.4000 ;
      RECT 15.0500 114.7000 15.5500 115.4000 ;
      RECT 14.2500 114.7000 14.7500 115.4000 ;
      RECT 13.4500 114.7000 13.9500 115.4000 ;
      RECT 12.6500 114.7000 13.1500 115.4000 ;
      RECT 11.8500 114.7000 12.3500 115.4000 ;
      RECT 11.0500 114.7000 11.5500 115.4000 ;
      RECT 10.2500 114.7000 10.7500 115.4000 ;
      RECT 0.0000 114.7000 9.9500 115.4000 ;
      RECT 0.0000 0.7000 118.4000 114.7000 ;
      RECT 111.8500 0.0000 118.4000 0.7000 ;
      RECT 111.0500 0.0000 111.5500 0.7000 ;
      RECT 110.2500 0.0000 110.7500 0.7000 ;
      RECT 109.4500 0.0000 109.9500 0.7000 ;
      RECT 108.6500 0.0000 109.1500 0.7000 ;
      RECT 107.8500 0.0000 108.3500 0.7000 ;
      RECT 107.0500 0.0000 107.5500 0.7000 ;
      RECT 106.2500 0.0000 106.7500 0.7000 ;
      RECT 105.4500 0.0000 105.9500 0.7000 ;
      RECT 104.6500 0.0000 105.1500 0.7000 ;
      RECT 103.8500 0.0000 104.3500 0.7000 ;
      RECT 103.0500 0.0000 103.5500 0.7000 ;
      RECT 102.2500 0.0000 102.7500 0.7000 ;
      RECT 101.4500 0.0000 101.9500 0.7000 ;
      RECT 100.6500 0.0000 101.1500 0.7000 ;
      RECT 99.8500 0.0000 100.3500 0.7000 ;
      RECT 99.0500 0.0000 99.5500 0.7000 ;
      RECT 98.2500 0.0000 98.7500 0.7000 ;
      RECT 97.4500 0.0000 97.9500 0.7000 ;
      RECT 96.6500 0.0000 97.1500 0.7000 ;
      RECT 95.8500 0.0000 96.3500 0.7000 ;
      RECT 95.0500 0.0000 95.5500 0.7000 ;
      RECT 94.2500 0.0000 94.7500 0.7000 ;
      RECT 93.4500 0.0000 93.9500 0.7000 ;
      RECT 92.6500 0.0000 93.1500 0.7000 ;
      RECT 91.8500 0.0000 92.3500 0.7000 ;
      RECT 91.0500 0.0000 91.5500 0.7000 ;
      RECT 90.2500 0.0000 90.7500 0.7000 ;
      RECT 89.4500 0.0000 89.9500 0.7000 ;
      RECT 88.6500 0.0000 89.1500 0.7000 ;
      RECT 87.8500 0.0000 88.3500 0.7000 ;
      RECT 87.0500 0.0000 87.5500 0.7000 ;
      RECT 86.2500 0.0000 86.7500 0.7000 ;
      RECT 85.4500 0.0000 85.9500 0.7000 ;
      RECT 84.6500 0.0000 85.1500 0.7000 ;
      RECT 83.8500 0.0000 84.3500 0.7000 ;
      RECT 83.0500 0.0000 83.5500 0.7000 ;
      RECT 82.2500 0.0000 82.7500 0.7000 ;
      RECT 81.4500 0.0000 81.9500 0.7000 ;
      RECT 80.6500 0.0000 81.1500 0.7000 ;
      RECT 79.8500 0.0000 80.3500 0.7000 ;
      RECT 79.0500 0.0000 79.5500 0.7000 ;
      RECT 78.2500 0.0000 78.7500 0.7000 ;
      RECT 77.4500 0.0000 77.9500 0.7000 ;
      RECT 76.6500 0.0000 77.1500 0.7000 ;
      RECT 75.8500 0.0000 76.3500 0.7000 ;
      RECT 75.0500 0.0000 75.5500 0.7000 ;
      RECT 74.2500 0.0000 74.7500 0.7000 ;
      RECT 73.4500 0.0000 73.9500 0.7000 ;
      RECT 72.6500 0.0000 73.1500 0.7000 ;
      RECT 71.8500 0.0000 72.3500 0.7000 ;
      RECT 71.0500 0.0000 71.5500 0.7000 ;
      RECT 70.2500 0.0000 70.7500 0.7000 ;
      RECT 69.4500 0.0000 69.9500 0.7000 ;
      RECT 68.6500 0.0000 69.1500 0.7000 ;
      RECT 67.8500 0.0000 68.3500 0.7000 ;
      RECT 67.0500 0.0000 67.5500 0.7000 ;
      RECT 66.2500 0.0000 66.7500 0.7000 ;
      RECT 65.4500 0.0000 65.9500 0.7000 ;
      RECT 64.6500 0.0000 65.1500 0.7000 ;
      RECT 63.8500 0.0000 64.3500 0.7000 ;
      RECT 63.0500 0.0000 63.5500 0.7000 ;
      RECT 62.2500 0.0000 62.7500 0.7000 ;
      RECT 61.4500 0.0000 61.9500 0.7000 ;
      RECT 60.6500 0.0000 61.1500 0.7000 ;
      RECT 59.8500 0.0000 60.3500 0.7000 ;
      RECT 59.0500 0.0000 59.5500 0.7000 ;
      RECT 58.2500 0.0000 58.7500 0.7000 ;
      RECT 57.4500 0.0000 57.9500 0.7000 ;
      RECT 56.6500 0.0000 57.1500 0.7000 ;
      RECT 55.8500 0.0000 56.3500 0.7000 ;
      RECT 55.0500 0.0000 55.5500 0.7000 ;
      RECT 54.2500 0.0000 54.7500 0.7000 ;
      RECT 53.4500 0.0000 53.9500 0.7000 ;
      RECT 52.6500 0.0000 53.1500 0.7000 ;
      RECT 51.8500 0.0000 52.3500 0.7000 ;
      RECT 51.0500 0.0000 51.5500 0.7000 ;
      RECT 50.2500 0.0000 50.7500 0.7000 ;
      RECT 49.4500 0.0000 49.9500 0.7000 ;
      RECT 48.6500 0.0000 49.1500 0.7000 ;
      RECT 47.8500 0.0000 48.3500 0.7000 ;
      RECT 47.0500 0.0000 47.5500 0.7000 ;
      RECT 46.2500 0.0000 46.7500 0.7000 ;
      RECT 45.4500 0.0000 45.9500 0.7000 ;
      RECT 44.6500 0.0000 45.1500 0.7000 ;
      RECT 43.8500 0.0000 44.3500 0.7000 ;
      RECT 43.0500 0.0000 43.5500 0.7000 ;
      RECT 42.2500 0.0000 42.7500 0.7000 ;
      RECT 41.4500 0.0000 41.9500 0.7000 ;
      RECT 40.6500 0.0000 41.1500 0.7000 ;
      RECT 39.8500 0.0000 40.3500 0.7000 ;
      RECT 39.0500 0.0000 39.5500 0.7000 ;
      RECT 38.2500 0.0000 38.7500 0.7000 ;
      RECT 37.4500 0.0000 37.9500 0.7000 ;
      RECT 36.6500 0.0000 37.1500 0.7000 ;
      RECT 35.8500 0.0000 36.3500 0.7000 ;
      RECT 35.0500 0.0000 35.5500 0.7000 ;
      RECT 34.2500 0.0000 34.7500 0.7000 ;
      RECT 33.4500 0.0000 33.9500 0.7000 ;
      RECT 32.6500 0.0000 33.1500 0.7000 ;
      RECT 31.8500 0.0000 32.3500 0.7000 ;
      RECT 31.0500 0.0000 31.5500 0.7000 ;
      RECT 30.2500 0.0000 30.7500 0.7000 ;
      RECT 29.4500 0.0000 29.9500 0.7000 ;
      RECT 28.6500 0.0000 29.1500 0.7000 ;
      RECT 27.8500 0.0000 28.3500 0.7000 ;
      RECT 27.0500 0.0000 27.5500 0.7000 ;
      RECT 26.2500 0.0000 26.7500 0.7000 ;
      RECT 25.4500 0.0000 25.9500 0.7000 ;
      RECT 24.6500 0.0000 25.1500 0.7000 ;
      RECT 23.8500 0.0000 24.3500 0.7000 ;
      RECT 23.0500 0.0000 23.5500 0.7000 ;
      RECT 22.2500 0.0000 22.7500 0.7000 ;
      RECT 21.4500 0.0000 21.9500 0.7000 ;
      RECT 20.6500 0.0000 21.1500 0.7000 ;
      RECT 19.8500 0.0000 20.3500 0.7000 ;
      RECT 19.0500 0.0000 19.5500 0.7000 ;
      RECT 18.2500 0.0000 18.7500 0.7000 ;
      RECT 17.4500 0.0000 17.9500 0.7000 ;
      RECT 16.6500 0.0000 17.1500 0.7000 ;
      RECT 15.8500 0.0000 16.3500 0.7000 ;
      RECT 15.0500 0.0000 15.5500 0.7000 ;
      RECT 14.2500 0.0000 14.7500 0.7000 ;
      RECT 13.4500 0.0000 13.9500 0.7000 ;
      RECT 12.6500 0.0000 13.1500 0.7000 ;
      RECT 11.8500 0.0000 12.3500 0.7000 ;
      RECT 11.0500 0.0000 11.5500 0.7000 ;
      RECT 10.2500 0.0000 10.7500 0.7000 ;
      RECT 0.0000 0.0000 9.9500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 69.7500 118.4000 115.4000 ;
      RECT 0.7000 69.4500 118.4000 69.7500 ;
      RECT 0.0000 65.7500 118.4000 69.4500 ;
      RECT 0.7000 65.4500 118.4000 65.7500 ;
      RECT 0.0000 61.7500 118.4000 65.4500 ;
      RECT 0.7000 61.4500 118.4000 61.7500 ;
      RECT 0.0000 57.7500 118.4000 61.4500 ;
      RECT 0.7000 57.4500 118.4000 57.7500 ;
      RECT 0.0000 53.7500 118.4000 57.4500 ;
      RECT 0.7000 53.4500 118.4000 53.7500 ;
      RECT 0.0000 49.7500 118.4000 53.4500 ;
      RECT 0.7000 49.4500 118.4000 49.7500 ;
      RECT 0.0000 45.7500 118.4000 49.4500 ;
      RECT 0.7000 45.4500 118.4000 45.7500 ;
      RECT 0.0000 0.0000 118.4000 45.4500 ;
    LAYER M4 ;
      RECT 0.0000 114.7250 118.4000 115.4000 ;
      RECT 8.1600 114.5600 113.8400 114.7250 ;
      RECT 0.0000 114.5600 6.8400 114.7250 ;
      RECT 115.1600 0.8400 118.4000 114.7250 ;
      RECT 113.1600 0.8400 113.8400 114.5600 ;
      RECT 8.1600 0.8400 111.8400 114.5600 ;
      RECT 6.1600 0.8400 6.8400 114.5600 ;
      RECT 113.1600 0.6750 118.4000 0.8400 ;
      RECT 6.1600 0.6750 111.8400 0.8400 ;
      RECT 0.0000 0.6750 4.8400 114.5600 ;
      RECT 0.0000 0.0000 118.4000 0.6750 ;
  END
END sram_w16

END LIBRARY
