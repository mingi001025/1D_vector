##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Tue Mar 11 14:00:38 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 458.0000 BY 455.6000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 181.9500 0.6000 182.0500 ;
    END
  END clk
  PIN sum_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.6500 0.0000 228.7500 0.6000 ;
    END
  END sum_out[159]
  PIN sum_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 227.6500 0.0000 227.7500 0.6000 ;
    END
  END sum_out[158]
  PIN sum_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.6500 0.0000 226.7500 0.6000 ;
    END
  END sum_out[157]
  PIN sum_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 225.6500 0.0000 225.7500 0.6000 ;
    END
  END sum_out[156]
  PIN sum_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 224.6500 0.0000 224.7500 0.6000 ;
    END
  END sum_out[155]
  PIN sum_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.6500 0.0000 223.7500 0.6000 ;
    END
  END sum_out[154]
  PIN sum_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 222.6500 0.0000 222.7500 0.6000 ;
    END
  END sum_out[153]
  PIN sum_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.6500 0.0000 221.7500 0.6000 ;
    END
  END sum_out[152]
  PIN sum_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 220.6500 0.0000 220.7500 0.6000 ;
    END
  END sum_out[151]
  PIN sum_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 219.6500 0.0000 219.7500 0.6000 ;
    END
  END sum_out[150]
  PIN sum_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 218.6500 0.0000 218.7500 0.6000 ;
    END
  END sum_out[149]
  PIN sum_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 217.6500 0.0000 217.7500 0.6000 ;
    END
  END sum_out[148]
  PIN sum_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 216.6500 0.0000 216.7500 0.6000 ;
    END
  END sum_out[147]
  PIN sum_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 215.6500 0.0000 215.7500 0.6000 ;
    END
  END sum_out[146]
  PIN sum_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 214.6500 0.0000 214.7500 0.6000 ;
    END
  END sum_out[145]
  PIN sum_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 213.6500 0.0000 213.7500 0.6000 ;
    END
  END sum_out[144]
  PIN sum_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 212.6500 0.0000 212.7500 0.6000 ;
    END
  END sum_out[143]
  PIN sum_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 211.6500 0.0000 211.7500 0.6000 ;
    END
  END sum_out[142]
  PIN sum_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 210.6500 0.0000 210.7500 0.6000 ;
    END
  END sum_out[141]
  PIN sum_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.6500 0.0000 209.7500 0.6000 ;
    END
  END sum_out[140]
  PIN sum_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 208.6500 0.0000 208.7500 0.6000 ;
    END
  END sum_out[139]
  PIN sum_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.6500 0.0000 207.7500 0.6000 ;
    END
  END sum_out[138]
  PIN sum_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 206.6500 0.0000 206.7500 0.6000 ;
    END
  END sum_out[137]
  PIN sum_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 205.6500 0.0000 205.7500 0.6000 ;
    END
  END sum_out[136]
  PIN sum_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.6500 0.0000 204.7500 0.6000 ;
    END
  END sum_out[135]
  PIN sum_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 203.6500 0.0000 203.7500 0.6000 ;
    END
  END sum_out[134]
  PIN sum_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.6500 0.0000 202.7500 0.6000 ;
    END
  END sum_out[133]
  PIN sum_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 201.6500 0.0000 201.7500 0.6000 ;
    END
  END sum_out[132]
  PIN sum_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 200.6500 0.0000 200.7500 0.6000 ;
    END
  END sum_out[131]
  PIN sum_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.6500 0.0000 199.7500 0.6000 ;
    END
  END sum_out[130]
  PIN sum_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 198.6500 0.0000 198.7500 0.6000 ;
    END
  END sum_out[129]
  PIN sum_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.6500 0.0000 197.7500 0.6000 ;
    END
  END sum_out[128]
  PIN sum_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 196.6500 0.0000 196.7500 0.6000 ;
    END
  END sum_out[127]
  PIN sum_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 195.6500 0.0000 195.7500 0.6000 ;
    END
  END sum_out[126]
  PIN sum_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 194.6500 0.0000 194.7500 0.6000 ;
    END
  END sum_out[125]
  PIN sum_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 193.6500 0.0000 193.7500 0.6000 ;
    END
  END sum_out[124]
  PIN sum_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 192.6500 0.0000 192.7500 0.6000 ;
    END
  END sum_out[123]
  PIN sum_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 191.6500 0.0000 191.7500 0.6000 ;
    END
  END sum_out[122]
  PIN sum_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 190.6500 0.0000 190.7500 0.6000 ;
    END
  END sum_out[121]
  PIN sum_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 189.6500 0.0000 189.7500 0.6000 ;
    END
  END sum_out[120]
  PIN sum_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 188.6500 0.0000 188.7500 0.6000 ;
    END
  END sum_out[119]
  PIN sum_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 187.6500 0.0000 187.7500 0.6000 ;
    END
  END sum_out[118]
  PIN sum_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 186.6500 0.0000 186.7500 0.6000 ;
    END
  END sum_out[117]
  PIN sum_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.6500 0.0000 185.7500 0.6000 ;
    END
  END sum_out[116]
  PIN sum_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 184.6500 0.0000 184.7500 0.6000 ;
    END
  END sum_out[115]
  PIN sum_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.6500 0.0000 183.7500 0.6000 ;
    END
  END sum_out[114]
  PIN sum_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 182.6500 0.0000 182.7500 0.6000 ;
    END
  END sum_out[113]
  PIN sum_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 181.6500 0.0000 181.7500 0.6000 ;
    END
  END sum_out[112]
  PIN sum_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.6500 0.0000 180.7500 0.6000 ;
    END
  END sum_out[111]
  PIN sum_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 179.6500 0.0000 179.7500 0.6000 ;
    END
  END sum_out[110]
  PIN sum_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.6500 0.0000 178.7500 0.6000 ;
    END
  END sum_out[109]
  PIN sum_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 177.6500 0.0000 177.7500 0.6000 ;
    END
  END sum_out[108]
  PIN sum_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 176.6500 0.0000 176.7500 0.6000 ;
    END
  END sum_out[107]
  PIN sum_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.6500 0.0000 175.7500 0.6000 ;
    END
  END sum_out[106]
  PIN sum_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 174.6500 0.0000 174.7500 0.6000 ;
    END
  END sum_out[105]
  PIN sum_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.6500 0.0000 173.7500 0.6000 ;
    END
  END sum_out[104]
  PIN sum_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 172.6500 0.0000 172.7500 0.6000 ;
    END
  END sum_out[103]
  PIN sum_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.6500 0.0000 171.7500 0.6000 ;
    END
  END sum_out[102]
  PIN sum_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 170.6500 0.0000 170.7500 0.6000 ;
    END
  END sum_out[101]
  PIN sum_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 169.6500 0.0000 169.7500 0.6000 ;
    END
  END sum_out[100]
  PIN sum_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.6500 0.0000 168.7500 0.6000 ;
    END
  END sum_out[99]
  PIN sum_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 167.6500 0.0000 167.7500 0.6000 ;
    END
  END sum_out[98]
  PIN sum_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.6500 0.0000 166.7500 0.6000 ;
    END
  END sum_out[97]
  PIN sum_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 165.6500 0.0000 165.7500 0.6000 ;
    END
  END sum_out[96]
  PIN sum_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 164.6500 0.0000 164.7500 0.6000 ;
    END
  END sum_out[95]
  PIN sum_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.6500 0.0000 163.7500 0.6000 ;
    END
  END sum_out[94]
  PIN sum_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 162.6500 0.0000 162.7500 0.6000 ;
    END
  END sum_out[93]
  PIN sum_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.6500 0.0000 161.7500 0.6000 ;
    END
  END sum_out[92]
  PIN sum_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 160.6500 0.0000 160.7500 0.6000 ;
    END
  END sum_out[91]
  PIN sum_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.6500 0.0000 159.7500 0.6000 ;
    END
  END sum_out[90]
  PIN sum_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.6500 0.0000 158.7500 0.6000 ;
    END
  END sum_out[89]
  PIN sum_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 157.6500 0.0000 157.7500 0.6000 ;
    END
  END sum_out[88]
  PIN sum_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.6500 0.0000 156.7500 0.6000 ;
    END
  END sum_out[87]
  PIN sum_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 155.6500 0.0000 155.7500 0.6000 ;
    END
  END sum_out[86]
  PIN sum_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 154.6500 0.0000 154.7500 0.6000 ;
    END
  END sum_out[85]
  PIN sum_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 153.6500 0.0000 153.7500 0.6000 ;
    END
  END sum_out[84]
  PIN sum_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 152.6500 0.0000 152.7500 0.6000 ;
    END
  END sum_out[83]
  PIN sum_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 151.6500 0.0000 151.7500 0.6000 ;
    END
  END sum_out[82]
  PIN sum_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 150.6500 0.0000 150.7500 0.6000 ;
    END
  END sum_out[81]
  PIN sum_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 149.6500 0.0000 149.7500 0.6000 ;
    END
  END sum_out[80]
  PIN sum_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 148.6500 0.0000 148.7500 0.6000 ;
    END
  END sum_out[79]
  PIN sum_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 147.6500 0.0000 147.7500 0.6000 ;
    END
  END sum_out[78]
  PIN sum_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 146.6500 0.0000 146.7500 0.6000 ;
    END
  END sum_out[77]
  PIN sum_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 145.6500 0.0000 145.7500 0.6000 ;
    END
  END sum_out[76]
  PIN sum_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 144.6500 0.0000 144.7500 0.6000 ;
    END
  END sum_out[75]
  PIN sum_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 143.6500 0.0000 143.7500 0.6000 ;
    END
  END sum_out[74]
  PIN sum_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 142.6500 0.0000 142.7500 0.6000 ;
    END
  END sum_out[73]
  PIN sum_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 141.6500 0.0000 141.7500 0.6000 ;
    END
  END sum_out[72]
  PIN sum_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 140.6500 0.0000 140.7500 0.6000 ;
    END
  END sum_out[71]
  PIN sum_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 139.6500 0.0000 139.7500 0.6000 ;
    END
  END sum_out[70]
  PIN sum_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 138.6500 0.0000 138.7500 0.6000 ;
    END
  END sum_out[69]
  PIN sum_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 137.6500 0.0000 137.7500 0.6000 ;
    END
  END sum_out[68]
  PIN sum_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 136.6500 0.0000 136.7500 0.6000 ;
    END
  END sum_out[67]
  PIN sum_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 135.6500 0.0000 135.7500 0.6000 ;
    END
  END sum_out[66]
  PIN sum_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 134.6500 0.0000 134.7500 0.6000 ;
    END
  END sum_out[65]
  PIN sum_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 133.6500 0.0000 133.7500 0.6000 ;
    END
  END sum_out[64]
  PIN sum_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 132.6500 0.0000 132.7500 0.6000 ;
    END
  END sum_out[63]
  PIN sum_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 131.6500 0.0000 131.7500 0.6000 ;
    END
  END sum_out[62]
  PIN sum_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 130.6500 0.0000 130.7500 0.6000 ;
    END
  END sum_out[61]
  PIN sum_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 129.6500 0.0000 129.7500 0.6000 ;
    END
  END sum_out[60]
  PIN sum_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 128.6500 0.0000 128.7500 0.6000 ;
    END
  END sum_out[59]
  PIN sum_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 127.6500 0.0000 127.7500 0.6000 ;
    END
  END sum_out[58]
  PIN sum_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 126.6500 0.0000 126.7500 0.6000 ;
    END
  END sum_out[57]
  PIN sum_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 125.6500 0.0000 125.7500 0.6000 ;
    END
  END sum_out[56]
  PIN sum_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 124.6500 0.0000 124.7500 0.6000 ;
    END
  END sum_out[55]
  PIN sum_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 123.6500 0.0000 123.7500 0.6000 ;
    END
  END sum_out[54]
  PIN sum_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 122.6500 0.0000 122.7500 0.6000 ;
    END
  END sum_out[53]
  PIN sum_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 121.6500 0.0000 121.7500 0.6000 ;
    END
  END sum_out[52]
  PIN sum_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 120.6500 0.0000 120.7500 0.6000 ;
    END
  END sum_out[51]
  PIN sum_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 119.6500 0.0000 119.7500 0.6000 ;
    END
  END sum_out[50]
  PIN sum_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 118.6500 0.0000 118.7500 0.6000 ;
    END
  END sum_out[49]
  PIN sum_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 117.6500 0.0000 117.7500 0.6000 ;
    END
  END sum_out[48]
  PIN sum_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 116.6500 0.0000 116.7500 0.6000 ;
    END
  END sum_out[47]
  PIN sum_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 115.6500 0.0000 115.7500 0.6000 ;
    END
  END sum_out[46]
  PIN sum_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 114.6500 0.0000 114.7500 0.6000 ;
    END
  END sum_out[45]
  PIN sum_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 113.6500 0.0000 113.7500 0.6000 ;
    END
  END sum_out[44]
  PIN sum_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 112.6500 0.0000 112.7500 0.6000 ;
    END
  END sum_out[43]
  PIN sum_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 111.6500 0.0000 111.7500 0.6000 ;
    END
  END sum_out[42]
  PIN sum_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 110.6500 0.0000 110.7500 0.6000 ;
    END
  END sum_out[41]
  PIN sum_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 109.6500 0.0000 109.7500 0.6000 ;
    END
  END sum_out[40]
  PIN sum_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 108.6500 0.0000 108.7500 0.6000 ;
    END
  END sum_out[39]
  PIN sum_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 107.6500 0.0000 107.7500 0.6000 ;
    END
  END sum_out[38]
  PIN sum_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 106.6500 0.0000 106.7500 0.6000 ;
    END
  END sum_out[37]
  PIN sum_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 105.6500 0.0000 105.7500 0.6000 ;
    END
  END sum_out[36]
  PIN sum_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 104.6500 0.0000 104.7500 0.6000 ;
    END
  END sum_out[35]
  PIN sum_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 103.6500 0.0000 103.7500 0.6000 ;
    END
  END sum_out[34]
  PIN sum_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 102.6500 0.0000 102.7500 0.6000 ;
    END
  END sum_out[33]
  PIN sum_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 101.6500 0.0000 101.7500 0.6000 ;
    END
  END sum_out[32]
  PIN sum_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 100.6500 0.0000 100.7500 0.6000 ;
    END
  END sum_out[31]
  PIN sum_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 99.6500 0.0000 99.7500 0.6000 ;
    END
  END sum_out[30]
  PIN sum_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 98.6500 0.0000 98.7500 0.6000 ;
    END
  END sum_out[29]
  PIN sum_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 97.6500 0.0000 97.7500 0.6000 ;
    END
  END sum_out[28]
  PIN sum_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.6500 0.0000 96.7500 0.6000 ;
    END
  END sum_out[27]
  PIN sum_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 95.6500 0.0000 95.7500 0.6000 ;
    END
  END sum_out[26]
  PIN sum_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 94.6500 0.0000 94.7500 0.6000 ;
    END
  END sum_out[25]
  PIN sum_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 93.6500 0.0000 93.7500 0.6000 ;
    END
  END sum_out[24]
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 92.6500 0.0000 92.7500 0.6000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 91.6500 0.0000 91.7500 0.6000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.6500 0.0000 90.7500 0.6000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.6500 0.0000 89.7500 0.6000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.6500 0.0000 88.7500 0.6000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.6500 0.0000 87.7500 0.6000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.6500 0.0000 86.7500 0.6000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.6500 0.0000 85.7500 0.6000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.6500 0.0000 84.7500 0.6000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 83.6500 0.0000 83.7500 0.6000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.6500 0.0000 82.7500 0.6000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.6500 0.0000 81.7500 0.6000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.6500 0.0000 80.7500 0.6000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.6500 0.0000 79.7500 0.6000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 78.6500 0.0000 78.7500 0.6000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.6500 0.0000 77.7500 0.6000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.6500 0.0000 76.7500 0.6000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 75.6500 0.0000 75.7500 0.6000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.6500 0.0000 74.7500 0.6000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.6500 0.0000 73.7500 0.6000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 72.6500 0.0000 72.7500 0.6000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.6500 0.0000 71.7500 0.6000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.6500 0.0000 70.7500 0.6000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.6500 0.0000 69.7500 0.6000 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 309.9500 0.6000 310.0500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 307.9500 0.6000 308.0500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 305.9500 0.6000 306.0500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 303.9500 0.6000 304.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 301.9500 0.6000 302.0500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 299.9500 0.6000 300.0500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 297.9500 0.6000 298.0500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 295.9500 0.6000 296.0500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 293.9500 0.6000 294.0500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 291.9500 0.6000 292.0500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 289.9500 0.6000 290.0500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 287.9500 0.6000 288.0500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 285.9500 0.6000 286.0500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 283.9500 0.6000 284.0500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 281.9500 0.6000 282.0500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 279.9500 0.6000 280.0500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 277.9500 0.6000 278.0500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 275.9500 0.6000 276.0500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 273.9500 0.6000 274.0500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 271.9500 0.6000 272.0500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 269.9500 0.6000 270.0500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 267.9500 0.6000 268.0500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 265.9500 0.6000 266.0500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 263.9500 0.6000 264.0500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 261.9500 0.6000 262.0500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 259.9500 0.6000 260.0500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 257.9500 0.6000 258.0500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 255.9500 0.6000 256.0500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 253.9500 0.6000 254.0500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 251.9500 0.6000 252.0500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 249.9500 0.6000 250.0500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 247.9500 0.6000 248.0500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 245.9500 0.6000 246.0500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 243.9500 0.6000 244.0500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 241.9500 0.6000 242.0500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 239.9500 0.6000 240.0500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 237.9500 0.6000 238.0500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 235.9500 0.6000 236.0500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 233.9500 0.6000 234.0500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 231.9500 0.6000 232.0500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 229.9500 0.6000 230.0500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 227.9500 0.6000 228.0500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 225.9500 0.6000 226.0500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 223.9500 0.6000 224.0500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 221.9500 0.6000 222.0500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 219.9500 0.6000 220.0500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 217.9500 0.6000 218.0500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.9500 0.6000 216.0500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.9500 0.6000 214.0500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 211.9500 0.6000 212.0500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.9500 0.6000 210.0500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 207.9500 0.6000 208.0500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.9500 0.6000 206.0500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 203.9500 0.6000 204.0500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 201.9500 0.6000 202.0500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 199.9500 0.6000 200.0500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 197.9500 0.6000 198.0500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.9500 0.6000 196.0500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 193.9500 0.6000 194.0500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 191.9500 0.6000 192.0500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 189.9500 0.6000 190.0500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 187.9500 0.6000 188.0500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 185.9500 0.6000 186.0500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 183.9500 0.6000 184.0500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 388.6500 0.0000 388.7500 0.6000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 387.6500 0.0000 387.7500 0.6000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 386.6500 0.0000 386.7500 0.6000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 385.6500 0.0000 385.7500 0.6000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 384.6500 0.0000 384.7500 0.6000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 383.6500 0.0000 383.7500 0.6000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.6500 0.0000 382.7500 0.6000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 381.6500 0.0000 381.7500 0.6000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 380.6500 0.0000 380.7500 0.6000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 379.6500 0.0000 379.7500 0.6000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 378.6500 0.0000 378.7500 0.6000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.6500 0.0000 377.7500 0.6000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 376.6500 0.0000 376.7500 0.6000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.6500 0.0000 375.7500 0.6000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 374.6500 0.0000 374.7500 0.6000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 373.6500 0.0000 373.7500 0.6000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.6500 0.0000 372.7500 0.6000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 371.6500 0.0000 371.7500 0.6000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.6500 0.0000 370.7500 0.6000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 369.6500 0.0000 369.7500 0.6000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 368.6500 0.0000 368.7500 0.6000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.6500 0.0000 367.7500 0.6000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 366.6500 0.0000 366.7500 0.6000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.6500 0.0000 365.7500 0.6000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 364.6500 0.0000 364.7500 0.6000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.6500 0.0000 363.7500 0.6000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 362.6500 0.0000 362.7500 0.6000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 361.6500 0.0000 361.7500 0.6000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 360.6500 0.0000 360.7500 0.6000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 359.6500 0.0000 359.7500 0.6000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 358.6500 0.0000 358.7500 0.6000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 357.6500 0.0000 357.7500 0.6000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 356.6500 0.0000 356.7500 0.6000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 355.6500 0.0000 355.7500 0.6000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 354.6500 0.0000 354.7500 0.6000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.6500 0.0000 353.7500 0.6000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 352.6500 0.0000 352.7500 0.6000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.6500 0.0000 351.7500 0.6000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 350.6500 0.0000 350.7500 0.6000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 349.6500 0.0000 349.7500 0.6000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.6500 0.0000 348.7500 0.6000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 347.6500 0.0000 347.7500 0.6000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.6500 0.0000 346.7500 0.6000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 345.6500 0.0000 345.7500 0.6000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 344.6500 0.0000 344.7500 0.6000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.6500 0.0000 343.7500 0.6000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 342.6500 0.0000 342.7500 0.6000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.6500 0.0000 341.7500 0.6000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 340.6500 0.0000 340.7500 0.6000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.6500 0.0000 339.7500 0.6000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 338.6500 0.0000 338.7500 0.6000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 337.6500 0.0000 337.7500 0.6000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.6500 0.0000 336.7500 0.6000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 335.6500 0.0000 335.7500 0.6000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.6500 0.0000 334.7500 0.6000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 333.6500 0.0000 333.7500 0.6000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 332.6500 0.0000 332.7500 0.6000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.6500 0.0000 331.7500 0.6000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 330.6500 0.0000 330.7500 0.6000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.6500 0.0000 329.7500 0.6000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 328.6500 0.0000 328.7500 0.6000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.6500 0.0000 327.7500 0.6000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 326.6500 0.0000 326.7500 0.6000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 325.6500 0.0000 325.7500 0.6000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.6500 0.0000 324.7500 0.6000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 323.6500 0.0000 323.7500 0.6000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.6500 0.0000 322.7500 0.6000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 321.6500 0.0000 321.7500 0.6000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 320.6500 0.0000 320.7500 0.6000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.6500 0.0000 319.7500 0.6000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 318.6500 0.0000 318.7500 0.6000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.6500 0.0000 317.7500 0.6000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 316.6500 0.0000 316.7500 0.6000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.6500 0.0000 315.7500 0.6000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 314.6500 0.0000 314.7500 0.6000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 313.6500 0.0000 313.7500 0.6000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.6500 0.0000 312.7500 0.6000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 311.6500 0.0000 311.7500 0.6000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.6500 0.0000 310.7500 0.6000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 309.6500 0.0000 309.7500 0.6000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 308.6500 0.0000 308.7500 0.6000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.6500 0.0000 307.7500 0.6000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 306.6500 0.0000 306.7500 0.6000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.6500 0.0000 305.7500 0.6000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 304.6500 0.0000 304.7500 0.6000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.6500 0.0000 303.7500 0.6000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 302.6500 0.0000 302.7500 0.6000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 301.6500 0.0000 301.7500 0.6000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.6500 0.0000 300.7500 0.6000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 299.6500 0.0000 299.7500 0.6000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.6500 0.0000 298.7500 0.6000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 297.6500 0.0000 297.7500 0.6000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 296.6500 0.0000 296.7500 0.6000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.6500 0.0000 295.7500 0.6000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 294.6500 0.0000 294.7500 0.6000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.6500 0.0000 293.7500 0.6000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 292.6500 0.0000 292.7500 0.6000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.6500 0.0000 291.7500 0.6000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 290.6500 0.0000 290.7500 0.6000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 289.6500 0.0000 289.7500 0.6000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 288.6500 0.0000 288.7500 0.6000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 287.6500 0.0000 287.7500 0.6000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.6500 0.0000 286.7500 0.6000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 285.6500 0.0000 285.7500 0.6000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 284.6500 0.0000 284.7500 0.6000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.6500 0.0000 283.7500 0.6000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 282.6500 0.0000 282.7500 0.6000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.6500 0.0000 281.7500 0.6000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 280.6500 0.0000 280.7500 0.6000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.6500 0.0000 279.7500 0.6000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 278.6500 0.0000 278.7500 0.6000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 277.6500 0.0000 277.7500 0.6000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.6500 0.0000 276.7500 0.6000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 275.6500 0.0000 275.7500 0.6000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.6500 0.0000 274.7500 0.6000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 273.6500 0.0000 273.7500 0.6000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 272.6500 0.0000 272.7500 0.6000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.6500 0.0000 271.7500 0.6000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 270.6500 0.0000 270.7500 0.6000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 269.6500 0.0000 269.7500 0.6000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 268.6500 0.0000 268.7500 0.6000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 267.6500 0.0000 267.7500 0.6000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 266.6500 0.0000 266.7500 0.6000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 265.6500 0.0000 265.7500 0.6000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 264.6500 0.0000 264.7500 0.6000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 263.6500 0.0000 263.7500 0.6000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 262.6500 0.0000 262.7500 0.6000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 261.6500 0.0000 261.7500 0.6000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 260.6500 0.0000 260.7500 0.6000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 259.6500 0.0000 259.7500 0.6000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 258.6500 0.0000 258.7500 0.6000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 257.6500 0.0000 257.7500 0.6000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 256.6500 0.0000 256.7500 0.6000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.6500 0.0000 255.7500 0.6000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 254.6500 0.0000 254.7500 0.6000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 253.6500 0.0000 253.7500 0.6000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.6500 0.0000 252.7500 0.6000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 251.6500 0.0000 251.7500 0.6000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.6500 0.0000 250.7500 0.6000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 249.6500 0.0000 249.7500 0.6000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 248.6500 0.0000 248.7500 0.6000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.6500 0.0000 247.7500 0.6000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 246.6500 0.0000 246.7500 0.6000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.6500 0.0000 245.7500 0.6000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 244.6500 0.0000 244.7500 0.6000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 243.6500 0.0000 243.7500 0.6000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 242.6500 0.0000 242.7500 0.6000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 241.6500 0.0000 241.7500 0.6000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 240.6500 0.0000 240.7500 0.6000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 239.6500 0.0000 239.7500 0.6000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 238.6500 0.0000 238.7500 0.6000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 237.6500 0.0000 237.7500 0.6000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 236.6500 0.0000 236.7500 0.6000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 235.6500 0.0000 235.7500 0.6000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 234.6500 0.0000 234.7500 0.6000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.6500 0.0000 233.7500 0.6000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 232.6500 0.0000 232.7500 0.6000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.6500 0.0000 231.7500 0.6000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 230.6500 0.0000 230.7500 0.6000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 229.6500 0.0000 229.7500 0.6000 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 179.9500 0.6000 180.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 177.9500 0.6000 178.0500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 175.9500 0.6000 176.0500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 173.9500 0.6000 174.0500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 171.9500 0.6000 172.0500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 169.9500 0.6000 170.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 167.9500 0.6000 168.0500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 165.9500 0.6000 166.0500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 163.9500 0.6000 164.0500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 161.9500 0.6000 162.0500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 159.9500 0.6000 160.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 157.9500 0.6000 158.0500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 155.9500 0.6000 156.0500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 153.9500 0.6000 154.0500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 151.9500 0.6000 152.0500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 149.9500 0.6000 150.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 147.9500 0.6000 148.0500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 145.9500 0.6000 146.0500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
    LAYER M3 ;
      RECT 0.0000 310.1500 458.0000 455.6000 ;
      RECT 0.7000 309.8500 458.0000 310.1500 ;
      RECT 0.0000 308.1500 458.0000 309.8500 ;
      RECT 0.7000 307.8500 458.0000 308.1500 ;
      RECT 0.0000 306.1500 458.0000 307.8500 ;
      RECT 0.7000 305.8500 458.0000 306.1500 ;
      RECT 0.0000 304.1500 458.0000 305.8500 ;
      RECT 0.7000 303.8500 458.0000 304.1500 ;
      RECT 0.0000 302.1500 458.0000 303.8500 ;
      RECT 0.7000 301.8500 458.0000 302.1500 ;
      RECT 0.0000 300.1500 458.0000 301.8500 ;
      RECT 0.7000 299.8500 458.0000 300.1500 ;
      RECT 0.0000 298.1500 458.0000 299.8500 ;
      RECT 0.7000 297.8500 458.0000 298.1500 ;
      RECT 0.0000 296.1500 458.0000 297.8500 ;
      RECT 0.7000 295.8500 458.0000 296.1500 ;
      RECT 0.0000 294.1500 458.0000 295.8500 ;
      RECT 0.7000 293.8500 458.0000 294.1500 ;
      RECT 0.0000 292.1500 458.0000 293.8500 ;
      RECT 0.7000 291.8500 458.0000 292.1500 ;
      RECT 0.0000 290.1500 458.0000 291.8500 ;
      RECT 0.7000 289.8500 458.0000 290.1500 ;
      RECT 0.0000 288.1500 458.0000 289.8500 ;
      RECT 0.7000 287.8500 458.0000 288.1500 ;
      RECT 0.0000 286.1500 458.0000 287.8500 ;
      RECT 0.7000 285.8500 458.0000 286.1500 ;
      RECT 0.0000 284.1500 458.0000 285.8500 ;
      RECT 0.7000 283.8500 458.0000 284.1500 ;
      RECT 0.0000 282.1500 458.0000 283.8500 ;
      RECT 0.7000 281.8500 458.0000 282.1500 ;
      RECT 0.0000 280.1500 458.0000 281.8500 ;
      RECT 0.7000 279.8500 458.0000 280.1500 ;
      RECT 0.0000 278.1500 458.0000 279.8500 ;
      RECT 0.7000 277.8500 458.0000 278.1500 ;
      RECT 0.0000 276.1500 458.0000 277.8500 ;
      RECT 0.7000 275.8500 458.0000 276.1500 ;
      RECT 0.0000 274.1500 458.0000 275.8500 ;
      RECT 0.7000 273.8500 458.0000 274.1500 ;
      RECT 0.0000 272.1500 458.0000 273.8500 ;
      RECT 0.7000 271.8500 458.0000 272.1500 ;
      RECT 0.0000 270.1500 458.0000 271.8500 ;
      RECT 0.7000 269.8500 458.0000 270.1500 ;
      RECT 0.0000 268.1500 458.0000 269.8500 ;
      RECT 0.7000 267.8500 458.0000 268.1500 ;
      RECT 0.0000 266.1500 458.0000 267.8500 ;
      RECT 0.7000 265.8500 458.0000 266.1500 ;
      RECT 0.0000 264.1500 458.0000 265.8500 ;
      RECT 0.7000 263.8500 458.0000 264.1500 ;
      RECT 0.0000 262.1500 458.0000 263.8500 ;
      RECT 0.7000 261.8500 458.0000 262.1500 ;
      RECT 0.0000 260.1500 458.0000 261.8500 ;
      RECT 0.7000 259.8500 458.0000 260.1500 ;
      RECT 0.0000 258.1500 458.0000 259.8500 ;
      RECT 0.7000 257.8500 458.0000 258.1500 ;
      RECT 0.0000 256.1500 458.0000 257.8500 ;
      RECT 0.7000 255.8500 458.0000 256.1500 ;
      RECT 0.0000 254.1500 458.0000 255.8500 ;
      RECT 0.7000 253.8500 458.0000 254.1500 ;
      RECT 0.0000 252.1500 458.0000 253.8500 ;
      RECT 0.7000 251.8500 458.0000 252.1500 ;
      RECT 0.0000 250.1500 458.0000 251.8500 ;
      RECT 0.7000 249.8500 458.0000 250.1500 ;
      RECT 0.0000 248.1500 458.0000 249.8500 ;
      RECT 0.7000 247.8500 458.0000 248.1500 ;
      RECT 0.0000 246.1500 458.0000 247.8500 ;
      RECT 0.7000 245.8500 458.0000 246.1500 ;
      RECT 0.0000 244.1500 458.0000 245.8500 ;
      RECT 0.7000 243.8500 458.0000 244.1500 ;
      RECT 0.0000 242.1500 458.0000 243.8500 ;
      RECT 0.7000 241.8500 458.0000 242.1500 ;
      RECT 0.0000 240.1500 458.0000 241.8500 ;
      RECT 0.7000 239.8500 458.0000 240.1500 ;
      RECT 0.0000 238.1500 458.0000 239.8500 ;
      RECT 0.7000 237.8500 458.0000 238.1500 ;
      RECT 0.0000 236.1500 458.0000 237.8500 ;
      RECT 0.7000 235.8500 458.0000 236.1500 ;
      RECT 0.0000 234.1500 458.0000 235.8500 ;
      RECT 0.7000 233.8500 458.0000 234.1500 ;
      RECT 0.0000 232.1500 458.0000 233.8500 ;
      RECT 0.7000 231.8500 458.0000 232.1500 ;
      RECT 0.0000 230.1500 458.0000 231.8500 ;
      RECT 0.7000 229.8500 458.0000 230.1500 ;
      RECT 0.0000 228.1500 458.0000 229.8500 ;
      RECT 0.7000 227.8500 458.0000 228.1500 ;
      RECT 0.0000 226.1500 458.0000 227.8500 ;
      RECT 0.7000 225.8500 458.0000 226.1500 ;
      RECT 0.0000 224.1500 458.0000 225.8500 ;
      RECT 0.7000 223.8500 458.0000 224.1500 ;
      RECT 0.0000 222.1500 458.0000 223.8500 ;
      RECT 0.7000 221.8500 458.0000 222.1500 ;
      RECT 0.0000 220.1500 458.0000 221.8500 ;
      RECT 0.7000 219.8500 458.0000 220.1500 ;
      RECT 0.0000 218.1500 458.0000 219.8500 ;
      RECT 0.7000 217.8500 458.0000 218.1500 ;
      RECT 0.0000 216.1500 458.0000 217.8500 ;
      RECT 0.7000 215.8500 458.0000 216.1500 ;
      RECT 0.0000 214.1500 458.0000 215.8500 ;
      RECT 0.7000 213.8500 458.0000 214.1500 ;
      RECT 0.0000 212.1500 458.0000 213.8500 ;
      RECT 0.7000 211.8500 458.0000 212.1500 ;
      RECT 0.0000 210.1500 458.0000 211.8500 ;
      RECT 0.7000 209.8500 458.0000 210.1500 ;
      RECT 0.0000 208.1500 458.0000 209.8500 ;
      RECT 0.7000 207.8500 458.0000 208.1500 ;
      RECT 0.0000 206.1500 458.0000 207.8500 ;
      RECT 0.7000 205.8500 458.0000 206.1500 ;
      RECT 0.0000 204.1500 458.0000 205.8500 ;
      RECT 0.7000 203.8500 458.0000 204.1500 ;
      RECT 0.0000 202.1500 458.0000 203.8500 ;
      RECT 0.7000 201.8500 458.0000 202.1500 ;
      RECT 0.0000 200.1500 458.0000 201.8500 ;
      RECT 0.7000 199.8500 458.0000 200.1500 ;
      RECT 0.0000 198.1500 458.0000 199.8500 ;
      RECT 0.7000 197.8500 458.0000 198.1500 ;
      RECT 0.0000 196.1500 458.0000 197.8500 ;
      RECT 0.7000 195.8500 458.0000 196.1500 ;
      RECT 0.0000 194.1500 458.0000 195.8500 ;
      RECT 0.7000 193.8500 458.0000 194.1500 ;
      RECT 0.0000 192.1500 458.0000 193.8500 ;
      RECT 0.7000 191.8500 458.0000 192.1500 ;
      RECT 0.0000 190.1500 458.0000 191.8500 ;
      RECT 0.7000 189.8500 458.0000 190.1500 ;
      RECT 0.0000 188.1500 458.0000 189.8500 ;
      RECT 0.7000 187.8500 458.0000 188.1500 ;
      RECT 0.0000 186.1500 458.0000 187.8500 ;
      RECT 0.7000 185.8500 458.0000 186.1500 ;
      RECT 0.0000 184.1500 458.0000 185.8500 ;
      RECT 0.7000 183.8500 458.0000 184.1500 ;
      RECT 0.0000 182.1500 458.0000 183.8500 ;
      RECT 0.7000 181.8500 458.0000 182.1500 ;
      RECT 0.0000 180.1500 458.0000 181.8500 ;
      RECT 0.7000 179.8500 458.0000 180.1500 ;
      RECT 0.0000 178.1500 458.0000 179.8500 ;
      RECT 0.7000 177.8500 458.0000 178.1500 ;
      RECT 0.0000 176.1500 458.0000 177.8500 ;
      RECT 0.7000 175.8500 458.0000 176.1500 ;
      RECT 0.0000 174.1500 458.0000 175.8500 ;
      RECT 0.7000 173.8500 458.0000 174.1500 ;
      RECT 0.0000 172.1500 458.0000 173.8500 ;
      RECT 0.7000 171.8500 458.0000 172.1500 ;
      RECT 0.0000 170.1500 458.0000 171.8500 ;
      RECT 0.7000 169.8500 458.0000 170.1500 ;
      RECT 0.0000 168.1500 458.0000 169.8500 ;
      RECT 0.7000 167.8500 458.0000 168.1500 ;
      RECT 0.0000 166.1500 458.0000 167.8500 ;
      RECT 0.7000 165.8500 458.0000 166.1500 ;
      RECT 0.0000 164.1500 458.0000 165.8500 ;
      RECT 0.7000 163.8500 458.0000 164.1500 ;
      RECT 0.0000 162.1500 458.0000 163.8500 ;
      RECT 0.7000 161.8500 458.0000 162.1500 ;
      RECT 0.0000 160.1500 458.0000 161.8500 ;
      RECT 0.7000 159.8500 458.0000 160.1500 ;
      RECT 0.0000 158.1500 458.0000 159.8500 ;
      RECT 0.7000 157.8500 458.0000 158.1500 ;
      RECT 0.0000 156.1500 458.0000 157.8500 ;
      RECT 0.7000 155.8500 458.0000 156.1500 ;
      RECT 0.0000 154.1500 458.0000 155.8500 ;
      RECT 0.7000 153.8500 458.0000 154.1500 ;
      RECT 0.0000 152.1500 458.0000 153.8500 ;
      RECT 0.7000 151.8500 458.0000 152.1500 ;
      RECT 0.0000 150.1500 458.0000 151.8500 ;
      RECT 0.7000 149.8500 458.0000 150.1500 ;
      RECT 0.0000 148.1500 458.0000 149.8500 ;
      RECT 0.7000 147.8500 458.0000 148.1500 ;
      RECT 0.0000 146.1500 458.0000 147.8500 ;
      RECT 0.7000 145.8500 458.0000 146.1500 ;
      RECT 0.0000 0.7600 458.0000 145.8500 ;
      RECT 388.9100 0.0000 458.0000 0.7600 ;
      RECT 387.9100 0.0000 388.4900 0.7600 ;
      RECT 386.9100 0.0000 387.4900 0.7600 ;
      RECT 385.9100 0.0000 386.4900 0.7600 ;
      RECT 384.9100 0.0000 385.4900 0.7600 ;
      RECT 383.9100 0.0000 384.4900 0.7600 ;
      RECT 382.9100 0.0000 383.4900 0.7600 ;
      RECT 381.9100 0.0000 382.4900 0.7600 ;
      RECT 380.9100 0.0000 381.4900 0.7600 ;
      RECT 379.9100 0.0000 380.4900 0.7600 ;
      RECT 378.9100 0.0000 379.4900 0.7600 ;
      RECT 377.9100 0.0000 378.4900 0.7600 ;
      RECT 376.9100 0.0000 377.4900 0.7600 ;
      RECT 375.9100 0.0000 376.4900 0.7600 ;
      RECT 374.9100 0.0000 375.4900 0.7600 ;
      RECT 373.9100 0.0000 374.4900 0.7600 ;
      RECT 372.9100 0.0000 373.4900 0.7600 ;
      RECT 371.9100 0.0000 372.4900 0.7600 ;
      RECT 370.9100 0.0000 371.4900 0.7600 ;
      RECT 369.9100 0.0000 370.4900 0.7600 ;
      RECT 368.9100 0.0000 369.4900 0.7600 ;
      RECT 367.9100 0.0000 368.4900 0.7600 ;
      RECT 366.9100 0.0000 367.4900 0.7600 ;
      RECT 365.9100 0.0000 366.4900 0.7600 ;
      RECT 364.9100 0.0000 365.4900 0.7600 ;
      RECT 363.9100 0.0000 364.4900 0.7600 ;
      RECT 362.9100 0.0000 363.4900 0.7600 ;
      RECT 361.9100 0.0000 362.4900 0.7600 ;
      RECT 360.9100 0.0000 361.4900 0.7600 ;
      RECT 359.9100 0.0000 360.4900 0.7600 ;
      RECT 358.9100 0.0000 359.4900 0.7600 ;
      RECT 357.9100 0.0000 358.4900 0.7600 ;
      RECT 356.9100 0.0000 357.4900 0.7600 ;
      RECT 355.9100 0.0000 356.4900 0.7600 ;
      RECT 354.9100 0.0000 355.4900 0.7600 ;
      RECT 353.9100 0.0000 354.4900 0.7600 ;
      RECT 352.9100 0.0000 353.4900 0.7600 ;
      RECT 351.9100 0.0000 352.4900 0.7600 ;
      RECT 350.9100 0.0000 351.4900 0.7600 ;
      RECT 349.9100 0.0000 350.4900 0.7600 ;
      RECT 348.9100 0.0000 349.4900 0.7600 ;
      RECT 347.9100 0.0000 348.4900 0.7600 ;
      RECT 346.9100 0.0000 347.4900 0.7600 ;
      RECT 345.9100 0.0000 346.4900 0.7600 ;
      RECT 344.9100 0.0000 345.4900 0.7600 ;
      RECT 343.9100 0.0000 344.4900 0.7600 ;
      RECT 342.9100 0.0000 343.4900 0.7600 ;
      RECT 341.9100 0.0000 342.4900 0.7600 ;
      RECT 340.9100 0.0000 341.4900 0.7600 ;
      RECT 339.9100 0.0000 340.4900 0.7600 ;
      RECT 338.9100 0.0000 339.4900 0.7600 ;
      RECT 337.9100 0.0000 338.4900 0.7600 ;
      RECT 336.9100 0.0000 337.4900 0.7600 ;
      RECT 335.9100 0.0000 336.4900 0.7600 ;
      RECT 334.9100 0.0000 335.4900 0.7600 ;
      RECT 333.9100 0.0000 334.4900 0.7600 ;
      RECT 332.9100 0.0000 333.4900 0.7600 ;
      RECT 331.9100 0.0000 332.4900 0.7600 ;
      RECT 330.9100 0.0000 331.4900 0.7600 ;
      RECT 329.9100 0.0000 330.4900 0.7600 ;
      RECT 328.9100 0.0000 329.4900 0.7600 ;
      RECT 327.9100 0.0000 328.4900 0.7600 ;
      RECT 326.9100 0.0000 327.4900 0.7600 ;
      RECT 325.9100 0.0000 326.4900 0.7600 ;
      RECT 324.9100 0.0000 325.4900 0.7600 ;
      RECT 323.9100 0.0000 324.4900 0.7600 ;
      RECT 322.9100 0.0000 323.4900 0.7600 ;
      RECT 321.9100 0.0000 322.4900 0.7600 ;
      RECT 320.9100 0.0000 321.4900 0.7600 ;
      RECT 319.9100 0.0000 320.4900 0.7600 ;
      RECT 318.9100 0.0000 319.4900 0.7600 ;
      RECT 317.9100 0.0000 318.4900 0.7600 ;
      RECT 316.9100 0.0000 317.4900 0.7600 ;
      RECT 315.9100 0.0000 316.4900 0.7600 ;
      RECT 314.9100 0.0000 315.4900 0.7600 ;
      RECT 313.9100 0.0000 314.4900 0.7600 ;
      RECT 312.9100 0.0000 313.4900 0.7600 ;
      RECT 311.9100 0.0000 312.4900 0.7600 ;
      RECT 310.9100 0.0000 311.4900 0.7600 ;
      RECT 309.9100 0.0000 310.4900 0.7600 ;
      RECT 308.9100 0.0000 309.4900 0.7600 ;
      RECT 307.9100 0.0000 308.4900 0.7600 ;
      RECT 306.9100 0.0000 307.4900 0.7600 ;
      RECT 305.9100 0.0000 306.4900 0.7600 ;
      RECT 304.9100 0.0000 305.4900 0.7600 ;
      RECT 303.9100 0.0000 304.4900 0.7600 ;
      RECT 302.9100 0.0000 303.4900 0.7600 ;
      RECT 301.9100 0.0000 302.4900 0.7600 ;
      RECT 300.9100 0.0000 301.4900 0.7600 ;
      RECT 299.9100 0.0000 300.4900 0.7600 ;
      RECT 298.9100 0.0000 299.4900 0.7600 ;
      RECT 297.9100 0.0000 298.4900 0.7600 ;
      RECT 296.9100 0.0000 297.4900 0.7600 ;
      RECT 295.9100 0.0000 296.4900 0.7600 ;
      RECT 294.9100 0.0000 295.4900 0.7600 ;
      RECT 293.9100 0.0000 294.4900 0.7600 ;
      RECT 292.9100 0.0000 293.4900 0.7600 ;
      RECT 291.9100 0.0000 292.4900 0.7600 ;
      RECT 290.9100 0.0000 291.4900 0.7600 ;
      RECT 289.9100 0.0000 290.4900 0.7600 ;
      RECT 288.9100 0.0000 289.4900 0.7600 ;
      RECT 287.9100 0.0000 288.4900 0.7600 ;
      RECT 286.9100 0.0000 287.4900 0.7600 ;
      RECT 285.9100 0.0000 286.4900 0.7600 ;
      RECT 284.9100 0.0000 285.4900 0.7600 ;
      RECT 283.9100 0.0000 284.4900 0.7600 ;
      RECT 282.9100 0.0000 283.4900 0.7600 ;
      RECT 281.9100 0.0000 282.4900 0.7600 ;
      RECT 280.9100 0.0000 281.4900 0.7600 ;
      RECT 279.9100 0.0000 280.4900 0.7600 ;
      RECT 278.9100 0.0000 279.4900 0.7600 ;
      RECT 277.9100 0.0000 278.4900 0.7600 ;
      RECT 276.9100 0.0000 277.4900 0.7600 ;
      RECT 275.9100 0.0000 276.4900 0.7600 ;
      RECT 274.9100 0.0000 275.4900 0.7600 ;
      RECT 273.9100 0.0000 274.4900 0.7600 ;
      RECT 272.9100 0.0000 273.4900 0.7600 ;
      RECT 271.9100 0.0000 272.4900 0.7600 ;
      RECT 270.9100 0.0000 271.4900 0.7600 ;
      RECT 269.9100 0.0000 270.4900 0.7600 ;
      RECT 268.9100 0.0000 269.4900 0.7600 ;
      RECT 267.9100 0.0000 268.4900 0.7600 ;
      RECT 266.9100 0.0000 267.4900 0.7600 ;
      RECT 265.9100 0.0000 266.4900 0.7600 ;
      RECT 264.9100 0.0000 265.4900 0.7600 ;
      RECT 263.9100 0.0000 264.4900 0.7600 ;
      RECT 262.9100 0.0000 263.4900 0.7600 ;
      RECT 261.9100 0.0000 262.4900 0.7600 ;
      RECT 260.9100 0.0000 261.4900 0.7600 ;
      RECT 259.9100 0.0000 260.4900 0.7600 ;
      RECT 258.9100 0.0000 259.4900 0.7600 ;
      RECT 257.9100 0.0000 258.4900 0.7600 ;
      RECT 256.9100 0.0000 257.4900 0.7600 ;
      RECT 255.9100 0.0000 256.4900 0.7600 ;
      RECT 254.9100 0.0000 255.4900 0.7600 ;
      RECT 253.9100 0.0000 254.4900 0.7600 ;
      RECT 252.9100 0.0000 253.4900 0.7600 ;
      RECT 251.9100 0.0000 252.4900 0.7600 ;
      RECT 250.9100 0.0000 251.4900 0.7600 ;
      RECT 249.9100 0.0000 250.4900 0.7600 ;
      RECT 248.9100 0.0000 249.4900 0.7600 ;
      RECT 247.9100 0.0000 248.4900 0.7600 ;
      RECT 246.9100 0.0000 247.4900 0.7600 ;
      RECT 245.9100 0.0000 246.4900 0.7600 ;
      RECT 244.9100 0.0000 245.4900 0.7600 ;
      RECT 243.9100 0.0000 244.4900 0.7600 ;
      RECT 242.9100 0.0000 243.4900 0.7600 ;
      RECT 241.9100 0.0000 242.4900 0.7600 ;
      RECT 240.9100 0.0000 241.4900 0.7600 ;
      RECT 239.9100 0.0000 240.4900 0.7600 ;
      RECT 238.9100 0.0000 239.4900 0.7600 ;
      RECT 237.9100 0.0000 238.4900 0.7600 ;
      RECT 236.9100 0.0000 237.4900 0.7600 ;
      RECT 235.9100 0.0000 236.4900 0.7600 ;
      RECT 234.9100 0.0000 235.4900 0.7600 ;
      RECT 233.9100 0.0000 234.4900 0.7600 ;
      RECT 232.9100 0.0000 233.4900 0.7600 ;
      RECT 231.9100 0.0000 232.4900 0.7600 ;
      RECT 230.9100 0.0000 231.4900 0.7600 ;
      RECT 229.9100 0.0000 230.4900 0.7600 ;
      RECT 228.9100 0.0000 229.4900 0.7600 ;
      RECT 227.9100 0.0000 228.4900 0.7600 ;
      RECT 226.9100 0.0000 227.4900 0.7600 ;
      RECT 225.9100 0.0000 226.4900 0.7600 ;
      RECT 224.9100 0.0000 225.4900 0.7600 ;
      RECT 223.9100 0.0000 224.4900 0.7600 ;
      RECT 222.9100 0.0000 223.4900 0.7600 ;
      RECT 221.9100 0.0000 222.4900 0.7600 ;
      RECT 220.9100 0.0000 221.4900 0.7600 ;
      RECT 219.9100 0.0000 220.4900 0.7600 ;
      RECT 218.9100 0.0000 219.4900 0.7600 ;
      RECT 217.9100 0.0000 218.4900 0.7600 ;
      RECT 216.9100 0.0000 217.4900 0.7600 ;
      RECT 215.9100 0.0000 216.4900 0.7600 ;
      RECT 214.9100 0.0000 215.4900 0.7600 ;
      RECT 213.9100 0.0000 214.4900 0.7600 ;
      RECT 212.9100 0.0000 213.4900 0.7600 ;
      RECT 211.9100 0.0000 212.4900 0.7600 ;
      RECT 210.9100 0.0000 211.4900 0.7600 ;
      RECT 209.9100 0.0000 210.4900 0.7600 ;
      RECT 208.9100 0.0000 209.4900 0.7600 ;
      RECT 207.9100 0.0000 208.4900 0.7600 ;
      RECT 206.9100 0.0000 207.4900 0.7600 ;
      RECT 205.9100 0.0000 206.4900 0.7600 ;
      RECT 204.9100 0.0000 205.4900 0.7600 ;
      RECT 203.9100 0.0000 204.4900 0.7600 ;
      RECT 202.9100 0.0000 203.4900 0.7600 ;
      RECT 201.9100 0.0000 202.4900 0.7600 ;
      RECT 200.9100 0.0000 201.4900 0.7600 ;
      RECT 199.9100 0.0000 200.4900 0.7600 ;
      RECT 198.9100 0.0000 199.4900 0.7600 ;
      RECT 197.9100 0.0000 198.4900 0.7600 ;
      RECT 196.9100 0.0000 197.4900 0.7600 ;
      RECT 195.9100 0.0000 196.4900 0.7600 ;
      RECT 194.9100 0.0000 195.4900 0.7600 ;
      RECT 193.9100 0.0000 194.4900 0.7600 ;
      RECT 192.9100 0.0000 193.4900 0.7600 ;
      RECT 191.9100 0.0000 192.4900 0.7600 ;
      RECT 190.9100 0.0000 191.4900 0.7600 ;
      RECT 189.9100 0.0000 190.4900 0.7600 ;
      RECT 188.9100 0.0000 189.4900 0.7600 ;
      RECT 187.9100 0.0000 188.4900 0.7600 ;
      RECT 186.9100 0.0000 187.4900 0.7600 ;
      RECT 185.9100 0.0000 186.4900 0.7600 ;
      RECT 184.9100 0.0000 185.4900 0.7600 ;
      RECT 183.9100 0.0000 184.4900 0.7600 ;
      RECT 182.9100 0.0000 183.4900 0.7600 ;
      RECT 181.9100 0.0000 182.4900 0.7600 ;
      RECT 180.9100 0.0000 181.4900 0.7600 ;
      RECT 179.9100 0.0000 180.4900 0.7600 ;
      RECT 178.9100 0.0000 179.4900 0.7600 ;
      RECT 177.9100 0.0000 178.4900 0.7600 ;
      RECT 176.9100 0.0000 177.4900 0.7600 ;
      RECT 175.9100 0.0000 176.4900 0.7600 ;
      RECT 174.9100 0.0000 175.4900 0.7600 ;
      RECT 173.9100 0.0000 174.4900 0.7600 ;
      RECT 172.9100 0.0000 173.4900 0.7600 ;
      RECT 171.9100 0.0000 172.4900 0.7600 ;
      RECT 170.9100 0.0000 171.4900 0.7600 ;
      RECT 169.9100 0.0000 170.4900 0.7600 ;
      RECT 168.9100 0.0000 169.4900 0.7600 ;
      RECT 167.9100 0.0000 168.4900 0.7600 ;
      RECT 166.9100 0.0000 167.4900 0.7600 ;
      RECT 165.9100 0.0000 166.4900 0.7600 ;
      RECT 164.9100 0.0000 165.4900 0.7600 ;
      RECT 163.9100 0.0000 164.4900 0.7600 ;
      RECT 162.9100 0.0000 163.4900 0.7600 ;
      RECT 161.9100 0.0000 162.4900 0.7600 ;
      RECT 160.9100 0.0000 161.4900 0.7600 ;
      RECT 159.9100 0.0000 160.4900 0.7600 ;
      RECT 158.9100 0.0000 159.4900 0.7600 ;
      RECT 157.9100 0.0000 158.4900 0.7600 ;
      RECT 156.9100 0.0000 157.4900 0.7600 ;
      RECT 155.9100 0.0000 156.4900 0.7600 ;
      RECT 154.9100 0.0000 155.4900 0.7600 ;
      RECT 153.9100 0.0000 154.4900 0.7600 ;
      RECT 152.9100 0.0000 153.4900 0.7600 ;
      RECT 151.9100 0.0000 152.4900 0.7600 ;
      RECT 150.9100 0.0000 151.4900 0.7600 ;
      RECT 149.9100 0.0000 150.4900 0.7600 ;
      RECT 148.9100 0.0000 149.4900 0.7600 ;
      RECT 147.9100 0.0000 148.4900 0.7600 ;
      RECT 146.9100 0.0000 147.4900 0.7600 ;
      RECT 145.9100 0.0000 146.4900 0.7600 ;
      RECT 144.9100 0.0000 145.4900 0.7600 ;
      RECT 143.9100 0.0000 144.4900 0.7600 ;
      RECT 142.9100 0.0000 143.4900 0.7600 ;
      RECT 141.9100 0.0000 142.4900 0.7600 ;
      RECT 140.9100 0.0000 141.4900 0.7600 ;
      RECT 139.9100 0.0000 140.4900 0.7600 ;
      RECT 138.9100 0.0000 139.4900 0.7600 ;
      RECT 137.9100 0.0000 138.4900 0.7600 ;
      RECT 136.9100 0.0000 137.4900 0.7600 ;
      RECT 135.9100 0.0000 136.4900 0.7600 ;
      RECT 134.9100 0.0000 135.4900 0.7600 ;
      RECT 133.9100 0.0000 134.4900 0.7600 ;
      RECT 132.9100 0.0000 133.4900 0.7600 ;
      RECT 131.9100 0.0000 132.4900 0.7600 ;
      RECT 130.9100 0.0000 131.4900 0.7600 ;
      RECT 129.9100 0.0000 130.4900 0.7600 ;
      RECT 128.9100 0.0000 129.4900 0.7600 ;
      RECT 127.9100 0.0000 128.4900 0.7600 ;
      RECT 126.9100 0.0000 127.4900 0.7600 ;
      RECT 125.9100 0.0000 126.4900 0.7600 ;
      RECT 124.9100 0.0000 125.4900 0.7600 ;
      RECT 123.9100 0.0000 124.4900 0.7600 ;
      RECT 122.9100 0.0000 123.4900 0.7600 ;
      RECT 121.9100 0.0000 122.4900 0.7600 ;
      RECT 120.9100 0.0000 121.4900 0.7600 ;
      RECT 119.9100 0.0000 120.4900 0.7600 ;
      RECT 118.9100 0.0000 119.4900 0.7600 ;
      RECT 117.9100 0.0000 118.4900 0.7600 ;
      RECT 116.9100 0.0000 117.4900 0.7600 ;
      RECT 115.9100 0.0000 116.4900 0.7600 ;
      RECT 114.9100 0.0000 115.4900 0.7600 ;
      RECT 113.9100 0.0000 114.4900 0.7600 ;
      RECT 112.9100 0.0000 113.4900 0.7600 ;
      RECT 111.9100 0.0000 112.4900 0.7600 ;
      RECT 110.9100 0.0000 111.4900 0.7600 ;
      RECT 109.9100 0.0000 110.4900 0.7600 ;
      RECT 108.9100 0.0000 109.4900 0.7600 ;
      RECT 107.9100 0.0000 108.4900 0.7600 ;
      RECT 106.9100 0.0000 107.4900 0.7600 ;
      RECT 105.9100 0.0000 106.4900 0.7600 ;
      RECT 104.9100 0.0000 105.4900 0.7600 ;
      RECT 103.9100 0.0000 104.4900 0.7600 ;
      RECT 102.9100 0.0000 103.4900 0.7600 ;
      RECT 101.9100 0.0000 102.4900 0.7600 ;
      RECT 100.9100 0.0000 101.4900 0.7600 ;
      RECT 99.9100 0.0000 100.4900 0.7600 ;
      RECT 98.9100 0.0000 99.4900 0.7600 ;
      RECT 97.9100 0.0000 98.4900 0.7600 ;
      RECT 96.9100 0.0000 97.4900 0.7600 ;
      RECT 95.9100 0.0000 96.4900 0.7600 ;
      RECT 94.9100 0.0000 95.4900 0.7600 ;
      RECT 93.9100 0.0000 94.4900 0.7600 ;
      RECT 92.9100 0.0000 93.4900 0.7600 ;
      RECT 91.9100 0.0000 92.4900 0.7600 ;
      RECT 90.9100 0.0000 91.4900 0.7600 ;
      RECT 89.9100 0.0000 90.4900 0.7600 ;
      RECT 88.9100 0.0000 89.4900 0.7600 ;
      RECT 87.9100 0.0000 88.4900 0.7600 ;
      RECT 86.9100 0.0000 87.4900 0.7600 ;
      RECT 85.9100 0.0000 86.4900 0.7600 ;
      RECT 84.9100 0.0000 85.4900 0.7600 ;
      RECT 83.9100 0.0000 84.4900 0.7600 ;
      RECT 82.9100 0.0000 83.4900 0.7600 ;
      RECT 81.9100 0.0000 82.4900 0.7600 ;
      RECT 80.9100 0.0000 81.4900 0.7600 ;
      RECT 79.9100 0.0000 80.4900 0.7600 ;
      RECT 78.9100 0.0000 79.4900 0.7600 ;
      RECT 77.9100 0.0000 78.4900 0.7600 ;
      RECT 76.9100 0.0000 77.4900 0.7600 ;
      RECT 75.9100 0.0000 76.4900 0.7600 ;
      RECT 74.9100 0.0000 75.4900 0.7600 ;
      RECT 73.9100 0.0000 74.4900 0.7600 ;
      RECT 72.9100 0.0000 73.4900 0.7600 ;
      RECT 71.9100 0.0000 72.4900 0.7600 ;
      RECT 70.9100 0.0000 71.4900 0.7600 ;
      RECT 69.9100 0.0000 70.4900 0.7600 ;
      RECT 0.0000 0.0000 69.4900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 458.0000 455.6000 ;
  END
END core

END LIBRARY
